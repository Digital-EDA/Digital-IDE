module SimpleAdd_1(
    input [8:0] a, b,
    output [8:0] c
);

    assign c = a + b;
    
    
endmodule //SimpleAdd


