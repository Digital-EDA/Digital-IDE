//------------------------------------------------------------------------------
// The confidential and proprietary information contained in this file may
// only be used by a person authorised under and to the extent permitted
// by a subsisting licensing agreement from ARM Limited or its affiliates.
//
//            (C) COPYRIGHT 2017 ARM Limited or its affiliates.
//                ALL RIGHTS RESERVED
//
// This entire notice must be reproduced on all copies of this file
// and copies of this file may only be made by a person if such person is
// permitted to do so under the terms of a subsisting license agreement
// from ARM Limited or its affiliates.
//
//  Version and Release Control Information:
//
//  File Revision       : $Revision: $
//  File Date           : $Date: $
//
//  Release Information : development
//
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Cortex-M0 DesignStart processor logic level
//------------------------------------------------------------------------------

module cortexm0ds_logic
(FCLK, SCLK, HCLK, DCLK, PORESETn, DBGRESETn, HRESETn,
SWCLKTCK, nTRST, HADDR, HBURST, HMASTLOCK, HPROT, HSIZE, HTRANS, HWDATA,
HWRITE, HRDATA, HREADY, HRESP, HMASTER, CODENSEQ, CODEHINTDE, SPECHTRANS
, SWDITMS, TDI, SWDO, SWDOEN, TDO, nTDOEN, DBGRESTART, DBGRESTARTED,
EDBGRQ, HALTED, NMI, IRQ, TXEV, RXEV, LOCKUP, SYSRESETREQ, STCALIB,
STCLKEN, IRQLATENCY, ECOREVNUM, GATEHCLK, SLEEPING, SLEEPDEEP, WAKEUP,
WICSENSE, SLEEPHOLDREQn, SLEEPHOLDACKn, WICENREQ, WICENACK, CDBGPWRUPREQ
, CDBGPWRUPACK, SE, RSTBYPASS, vis_r0_o, vis_r1_o, vis_r2_o, vis_r3_o,
vis_r4_o, vis_r5_o, vis_r6_o, vis_r7_o, vis_r8_o, vis_r9_o, vis_r10_o,
vis_r11_o, vis_r12_o, vis_r14_o, vis_msp_o, vis_psp_o, vis_pc_o,
vis_apsr_o, vis_tbit_o, vis_ipsr_o, vis_control_o, vis_primask_o);

output [31:0] HADDR;
output [2:0] HBURST;
output [3:0] HPROT;
output [2:0] HSIZE;
output [1:0] HTRANS;
output [31:0] HWDATA;
input [31:0] HRDATA;
output [2:0] CODEHINTDE;
input [31:0] IRQ;
input [25:0] STCALIB;
input [7:0] IRQLATENCY;
input [27:0] ECOREVNUM;
output [33:0] WICSENSE;
output [31:0] vis_r0_o;
output [31:0] vis_r1_o;
output [31:0] vis_r2_o;
output [31:0] vis_r3_o;
output [31:0] vis_r4_o;
output [31:0] vis_r5_o;
output [31:0] vis_r6_o;
output [31:0] vis_r7_o;
output [31:0] vis_r8_o;
output [31:0] vis_r9_o;
output [31:0] vis_r10_o;
output [31:0] vis_r11_o;
output [31:0] vis_r12_o;
output [31:0] vis_r14_o;
output [29:0] vis_msp_o;
output [29:0] vis_psp_o;
output [30:0] vis_pc_o;
output [3:0] vis_apsr_o;
output [5:0] vis_ipsr_o;
input FCLK;
input SCLK;
input HCLK;
input DCLK;
input PORESETn;
input DBGRESETn;
input HRESETn;
input SWCLKTCK;
input nTRST;
input HREADY;
input HRESP;
input SWDITMS;
input TDI;
input DBGRESTART;
input EDBGRQ;
input NMI;
input RXEV;
input STCLKEN;
input SLEEPHOLDREQn;
input WICENREQ;
input CDBGPWRUPACK;
input SE;
input RSTBYPASS;
output HMASTLOCK;
output HWRITE;
output HMASTER;
output CODENSEQ;
output SPECHTRANS;
output SWDO;
output SWDOEN;
output TDO;
output nTDOEN;
output DBGRESTARTED;
output HALTED;
output TXEV;
output LOCKUP;
output SYSRESETREQ;
output GATEHCLK;
output SLEEPING;
output SLEEPDEEP;
output WAKEUP;
output SLEEPHOLDACKn;
output WICENACK;
output CDBGPWRUPREQ;
output vis_tbit_o;
output vis_control_o;
output vis_primask_o;

wire Fmdhu6, Qmdhu6, Pndhu6, Oodhu6, Npdhu6, Qqdhu6, Fsdhu6, Stdhu6, Fvdhu6, Qwdhu6;
wire Jydhu6, C0ehu6, S1ehu6, L3ehu6, E5ehu6, T6ehu6, L8ehu6, Caehu6, Qbehu6, Edehu6;
wire Seehu6, Ggehu6, Uhehu6, Ijehu6, Wkehu6, Kmehu6, Ynehu6, Mpehu6, Arehu6, Osehu6;
wire Cuehu6, Qvehu6, Exehu6, Syehu6, G0fhu6, U1fhu6, I3fhu6, W4fhu6, K6fhu6, Y7fhu6;
wire M9fhu6, Abfhu6, Ocfhu6, Cefhu6, Qffhu6, Dhfhu6, Qifhu6, Dkfhu6, Qlfhu6, Dnfhu6;
wire Qofhu6, Dqfhu6, Vrfhu6, Ntfhu6, Ivfhu6, Dxfhu6, Yyfhu6, R0ghu6, N2ghu6, H4ghu6;
wire H6ghu6, Y7ghu6, V9ghu6, Sbghu6, Ndghu6, Gfghu6, Ahghu6, Righu6, Ikghu6, Zlghu6;
wire Qnghu6, Npghu6, Krghu6, Ftghu6, Dvghu6, Bxghu6, Yyghu6, T0hhu6, H2hhu6, S3hhu6;
wire E5hhu6, R6hhu6, D8hhu6, P9hhu6, Hbhhu6, Vchhu6, Jehhu6, Aghhu6, Qhhhu6, Ijhhu6;
wire Alhhu6, Smhhu6, Kohhu6, Wphhu6, Drhhu6, Kshhu6, Rthhu6, Yuhhu6, Gwhhu6, Oxhhu6;
wire Wyhhu6, E0ihu6, M1ihu6, U2ihu6, C4ihu6, K5ihu6, S6ihu6, A8ihu6, I9ihu6, Qaihu6;
wire Ybihu6, Gdihu6, Oeihu6, Wfihu6, Ehihu6, Miihu6, Ujihu6, Clihu6, Kmihu6, Snihu6;
wire Apihu6, Iqihu6, Qrihu6, Ysihu6, Guihu6, Ovihu6, Wwihu6, Eyihu6, Mzihu6, U0jhu6;
wire C2jhu6, K3jhu6, S4jhu6, A6jhu6, I7jhu6, Q8jhu6, Y9jhu6, Gbjhu6, Ocjhu6, Wdjhu6;
wire Efjhu6, Mgjhu6, Uhjhu6, Cjjhu6, Kkjhu6, Sljhu6, Anjhu6, Iojhu6, Qpjhu6, Yqjhu6;
wire Gsjhu6, Otjhu6, Wujhu6, Ewjhu6, Mxjhu6, Uyjhu6, C0khu6, K1khu6, S2khu6, A4khu6;
wire I5khu6, Q6khu6, Y7khu6, G9khu6, Oakhu6, Wbkhu6, Edkhu6, Mekhu6, Ufkhu6, Chkhu6;
wire Kikhu6, Sjkhu6, Alkhu6, Imkhu6, Qnkhu6, Yokhu6, Gqkhu6, Orkhu6, Wskhu6, Eukhu6;
wire Mvkhu6, Uwkhu6, Cykhu6, Kzkhu6, S0lhu6, A2lhu6, I3lhu6, Q4lhu6, Y5lhu6, G7lhu6;
wire O8lhu6, W9lhu6, Eblhu6, Lclhu6, Sdlhu6, Zelhu6, Gglhu6, Nhlhu6, Uilhu6, Bklhu6;
wire Illhu6, Pmlhu6, Wnlhu6, Dplhu6, Kqlhu6, Rrlhu6, Yslhu6, Fulhu6, Mvlhu6, Twlhu6;
wire Aylhu6, Hzlhu6, O0mhu6, V1mhu6, C3mhu6, J4mhu6, Q5mhu6, X6mhu6, E8mhu6, L9mhu6;
wire Samhu6, Zbmhu6, Gdmhu6, Nemhu6, Ufmhu6, Bhmhu6, Iimhu6, Pjmhu6, Wkmhu6, Dmmhu6;
wire Knmhu6, Romhu6, Ypmhu6, Frmhu6, Msmhu6, Ttmhu6, Avmhu6, Hwmhu6, Vxmhu6, Jzmhu6;
wire R0nhu6, A2nhu6, N3nhu6, I5nhu6, B7nhu6, Q8nhu6, Fanhu6, Ubnhu6, Jdnhu6, Yenhu6;
wire Rgnhu6, Pinhu6, Hknhu6, Ulnhu6, Fnnhu6, Tonhu6, Iqnhu6, Rrnhu6, Dtnhu6, Punhu6;
wire Gwnhu6, Cynhu6, Lznhu6, X0ohu6, G2ohu6, S3ohu6, O5ohu6, Q7ohu6, M9ohu6, R9ohu6;
wire W9ohu6, Daohu6, Kaohu6, Raohu6, Yaohu6, Fbohu6, Mbohu6, Tbohu6, Acohu6, Hcohu6;
wire Ocohu6, Vcohu6, Cdohu6, Jdohu6, Qdohu6, Xdohu6, Eeohu6, Leohu6, Seohu6, Zeohu6;
wire Gfohu6, Nfohu6, Ufohu6, Bgohu6, Igohu6, Pgohu6, Wgohu6, Dhohu6, Khohu6, Rhohu6;
wire Yhohu6, Fiohu6, Miohu6, Tiohu6, Ajohu6, Hjohu6, Ojohu6, Vjohu6, Ckohu6, Jkohu6;
wire Qkohu6, Xkohu6, Elohu6, Llohu6, Slohu6, Zlohu6, Gmohu6, Nmohu6, Umohu6, Bnohu6;
wire Inohu6, Pnohu6, Wnohu6, Doohu6, Koohu6, Roohu6, Yoohu6, Fpohu6, Mpohu6, Tpohu6;
wire Aqohu6, Hqohu6, Oqohu6, Vqohu6, Crohu6, Jrohu6, Qrohu6, Xrohu6, Esohu6, Lsohu6;
wire Ssohu6, Zsohu6, Gtohu6, Ntohu6, Utohu6, Buohu6, Iuohu6, Puohu6, Wuohu6, Dvohu6;
wire Kvohu6, Rvohu6, Yvohu6, Fwohu6, Mwohu6, Twohu6, Axohu6, Hxohu6, Oxohu6, Vxohu6;
wire Cyohu6, Jyohu6, Qyohu6, Xyohu6, Ezohu6, Lzohu6, Szohu6, Zzohu6, G0phu6, N0phu6;
wire U0phu6, B1phu6, I1phu6, P1phu6, W1phu6, D2phu6, K2phu6, R2phu6, Y2phu6, F3phu6;
wire M3phu6, T3phu6, A4phu6, H4phu6, O4phu6, V4phu6, C5phu6, J5phu6, Q5phu6, X5phu6;
wire E6phu6, L6phu6, S6phu6, Z6phu6, G7phu6, N7phu6, U7phu6, B8phu6, I8phu6, P8phu6;
wire W8phu6, D9phu6, K9phu6, R9phu6, Y9phu6, Faphu6, Maphu6, Taphu6, Abphu6, Hbphu6;
wire Obphu6, Vbphu6, Ccphu6, Jcphu6, Qcphu6, Xcphu6, Edphu6, Ldphu6, Sdphu6, Zdphu6;
wire Gephu6, Nephu6, Uephu6, Bfphu6, Ifphu6, Pfphu6, Wfphu6, Dgphu6, Kgphu6, Rgphu6;
wire Ygphu6, Fhphu6, Mhphu6, Thphu6, Aiphu6, Hiphu6, Oiphu6, Viphu6, Cjphu6, Jjphu6;
wire Qjphu6, Xjphu6, Ekphu6, Lkphu6, Skphu6, Zkphu6, Glphu6, Nlphu6, Ulphu6, Bmphu6;
wire Imphu6, Pmphu6, Wmphu6, Dnphu6, Knphu6, Rnphu6, Ynphu6, Fophu6, Mophu6, Tophu6;
wire Apphu6, Hpphu6, Opphu6, Vpphu6, Cqphu6, Jqphu6, Qqphu6, Xqphu6, Erphu6, Lrphu6;
wire Srphu6, Zrphu6, Gsphu6, Nsphu6, Usphu6, Btphu6, Itphu6, Ptphu6, Wtphu6, Duphu6;
wire Kuphu6, Ruphu6, Yuphu6, Fvphu6, Mvphu6, Tvphu6, Awphu6, Hwphu6, Owphu6, Vwphu6;
wire Cxphu6, Jxphu6, Qxphu6, Xxphu6, Eyphu6, Lyphu6, Syphu6, Zyphu6, Gzphu6, Nzphu6;
wire Uzphu6, B0qhu6, I0qhu6, P0qhu6, W0qhu6, D1qhu6, K1qhu6, R1qhu6, Y1qhu6, F2qhu6;
wire M2qhu6, T2qhu6, A3qhu6, H3qhu6, O3qhu6, V3qhu6, C4qhu6, J4qhu6, Q4qhu6, X4qhu6;
wire E5qhu6, L5qhu6, S5qhu6, Z5qhu6, G6qhu6, N6qhu6, U6qhu6, B7qhu6, I7qhu6, P7qhu6;
wire W7qhu6, D8qhu6, K8qhu6, R8qhu6, Y8qhu6, F9qhu6, M9qhu6, T9qhu6, Aaqhu6, Haqhu6;
wire Oaqhu6, Vaqhu6, Cbqhu6, Jbqhu6, Qbqhu6, Xbqhu6, Ecqhu6, Lcqhu6, Scqhu6, Zcqhu6;
wire Gdqhu6, Ndqhu6, Udqhu6, Beqhu6, Ieqhu6, Peqhu6, Weqhu6, Dfqhu6, Kfqhu6, Rfqhu6;
wire Yfqhu6, Fgqhu6, Mgqhu6, Tgqhu6, Ahqhu6, Hhqhu6, Ohqhu6, Vhqhu6, Ciqhu6, Jiqhu6;
wire Qiqhu6, Xiqhu6, Ejqhu6, Ljqhu6, Sjqhu6, Zjqhu6, Gkqhu6, Nkqhu6, Ukqhu6, Blqhu6;
wire Ilqhu6, Plqhu6, Wlqhu6, Dmqhu6, Kmqhu6, Rmqhu6, Ymqhu6, Fnqhu6, Mnqhu6, Tnqhu6;
wire Aoqhu6, Hoqhu6, Ooqhu6, Voqhu6, Cpqhu6, Jpqhu6, Qpqhu6, Xpqhu6, Eqqhu6, Lqqhu6;
wire Sqqhu6, Zqqhu6, Grqhu6, Nrqhu6, Urqhu6, Bsqhu6, Isqhu6, Psqhu6, Wsqhu6, Dtqhu6;
wire Ktqhu6, Rtqhu6, Ytqhu6, Fuqhu6, Muqhu6, Tuqhu6, Avqhu6, Hvqhu6, Ovqhu6, Vvqhu6;
wire Cwqhu6, Jwqhu6, Qwqhu6, Xwqhu6, Exqhu6, Lxqhu6, Sxqhu6, Zxqhu6, Gyqhu6, Nyqhu6;
wire Uyqhu6, Bzqhu6, Izqhu6, Pzqhu6, Wzqhu6, D0rhu6, K0rhu6, R0rhu6, Y0rhu6, F1rhu6;
wire M1rhu6, T1rhu6, A2rhu6, H2rhu6, O2rhu6, V2rhu6, C3rhu6, J3rhu6, Q3rhu6, X3rhu6;
wire E4rhu6, L4rhu6, S4rhu6, Z4rhu6, G5rhu6, N5rhu6, U5rhu6, B6rhu6, I6rhu6, P6rhu6;
wire W6rhu6, D7rhu6, K7rhu6, R7rhu6, Y7rhu6, F8rhu6, M8rhu6, T8rhu6, A9rhu6, H9rhu6;
wire O9rhu6, V9rhu6, Carhu6, Jarhu6, Qarhu6, Xarhu6, Ebrhu6, Lbrhu6, Sbrhu6, Zbrhu6;
wire Gcrhu6, Ncrhu6, Ucrhu6, Bdrhu6, Idrhu6, Pdrhu6, Wdrhu6, Derhu6, Kerhu6, Rerhu6;
wire Yerhu6, Ffrhu6, Mfrhu6, Tfrhu6, Agrhu6, Hgrhu6, Ogrhu6, Vgrhu6, Chrhu6, Jhrhu6;
wire Qhrhu6, Xhrhu6, Eirhu6, Lirhu6, Sirhu6, Zirhu6, Gjrhu6, Njrhu6, Ujrhu6, Bkrhu6;
wire Ikrhu6, Pkrhu6, Wkrhu6, Dlrhu6, Klrhu6, Rlrhu6, Ylrhu6, Fmrhu6, Mmrhu6, Tmrhu6;
wire Anrhu6, Hnrhu6, Onrhu6, Vnrhu6, Corhu6, Jorhu6, Qorhu6, Xorhu6, Eprhu6, Lprhu6;
wire Sprhu6, Zprhu6, Gqrhu6, Nqrhu6, Uqrhu6, Brrhu6, Irrhu6, Prrhu6, Wrrhu6, Dsrhu6;
wire Ksrhu6, Rsrhu6, Ysrhu6, Ftrhu6, Mtrhu6, Ttrhu6, Aurhu6, Hurhu6, Ourhu6, Vurhu6;
wire Cvrhu6, Jvrhu6, Qvrhu6, Xvrhu6, Ewrhu6, Lwrhu6, Swrhu6, Zwrhu6, Gxrhu6, Nxrhu6;
wire Uxrhu6, Byrhu6, Iyrhu6, Pyrhu6, Wyrhu6, Dzrhu6, Kzrhu6, Rzrhu6, Yzrhu6, F0shu6;
wire M0shu6, T0shu6, A1shu6, H1shu6, O1shu6, V1shu6, C2shu6, J2shu6, Q2shu6, X2shu6;
wire E3shu6, L3shu6, S3shu6, Z3shu6, G4shu6, N4shu6, U4shu6, B5shu6, I5shu6, P5shu6;
wire W5shu6, D6shu6, K6shu6, R6shu6, Y6shu6, F7shu6, M7shu6, T7shu6, A8shu6, H8shu6;
wire O8shu6, V8shu6, C9shu6, J9shu6, Q9shu6, X9shu6, Eashu6, Lashu6, Sashu6, Zashu6;
wire Gbshu6, Nbshu6, Ubshu6, Bcshu6, Icshu6, Pcshu6, Wcshu6, Ddshu6, Kdshu6, Rdshu6;
wire Ydshu6, Feshu6, Meshu6, Teshu6, Afshu6, Hfshu6, Ofshu6, Vfshu6, Cgshu6, Jgshu6;
wire Qgshu6, Xgshu6, Ehshu6, Lhshu6, Shshu6, Zhshu6, Gishu6, Nishu6, Uishu6, Bjshu6;
wire Ijshu6, Pjshu6, Wjshu6, Dkshu6, Kkshu6, Rkshu6, Ykshu6, Flshu6, Mlshu6, Tlshu6;
wire Amshu6, Hmshu6, Omshu6, Vmshu6, Cnshu6, Jnshu6, Qnshu6, Xnshu6, Eoshu6, Loshu6;
wire Soshu6, Zoshu6, Gpshu6, Npshu6, Upshu6, Bqshu6, Iqshu6, Pqshu6, Wqshu6, Drshu6;
wire Krshu6, Rrshu6, Yrshu6, Fsshu6, Msshu6, Tsshu6, Atshu6, Htshu6, Otshu6, Vtshu6;
wire Cushu6, Jushu6, Qushu6, Xushu6, Evshu6, Lvshu6, Svshu6, Zvshu6, Gwshu6, Nwshu6;
wire Uwshu6, Bxshu6, Ixshu6, Pxshu6, Wxshu6, Dyshu6, Kyshu6, Ryshu6, Yyshu6, Fzshu6;
wire Mzshu6, Tzshu6, A0thu6, H0thu6, O0thu6, V0thu6, C1thu6, J1thu6, Q1thu6, X1thu6;
wire E2thu6, L2thu6, S2thu6, Z2thu6, G3thu6, N3thu6, U3thu6, B4thu6, I4thu6, P4thu6;
wire W4thu6, D5thu6, K5thu6, R5thu6, Y5thu6, F6thu6, M6thu6, T6thu6, A7thu6, H7thu6;
wire O7thu6, V7thu6, C8thu6, J8thu6, Q8thu6, X8thu6, E9thu6, L9thu6, S9thu6, Z9thu6;
wire Gathu6, Nathu6, Uathu6, Bbthu6, Ibthu6, Pbthu6, Wbthu6, Dcthu6, Kcthu6, Rcthu6;
wire Ycthu6, Fdthu6, Mdthu6, Tdthu6, Aethu6, Hethu6, Oethu6, Vethu6, Cfthu6, Jfthu6;
wire Qfthu6, Xfthu6, Egthu6, Lgthu6, Sgthu6, Zgthu6, Ghthu6, Nhthu6, Uhthu6, Bithu6;
wire Iithu6, Pithu6, Withu6, Djthu6, Kjthu6, Rjthu6, Yjthu6, Fkthu6, Mkthu6, Tkthu6;
wire Althu6, Hlthu6, Olthu6, Vlthu6, Cmthu6, Jmthu6, Qmthu6, Xmthu6, Enthu6, Lnthu6;
wire Snthu6, Znthu6, Gothu6, Nothu6, Uothu6, Bpthu6, Ipthu6, Ppthu6, Wpthu6, Dqthu6;
wire Kqthu6, Rqthu6, Yqthu6, Frthu6, Mrthu6, Trthu6, Asthu6, Hsthu6, Osthu6, Vsthu6;
wire Ctthu6, Jtthu6, Qtthu6, Xtthu6, Euthu6, Luthu6, Suthu6, Zuthu6, Gvthu6, Nvthu6;
wire Uvthu6, Bwthu6, Iwthu6, Pwthu6, Wwthu6, Dxthu6, Kxthu6, Rxthu6, Yxthu6, Fythu6;
wire Mythu6, Tythu6, Azthu6, Hzthu6, Ozthu6, Vzthu6, C0uhu6, J0uhu6, Q0uhu6, X0uhu6;
wire E1uhu6, L1uhu6, S1uhu6, Z1uhu6, G2uhu6, N2uhu6, U2uhu6, B3uhu6, I3uhu6, P3uhu6;
wire W3uhu6, D4uhu6, K4uhu6, R4uhu6, Y4uhu6, F5uhu6, M5uhu6, T5uhu6, A6uhu6, H6uhu6;
wire O6uhu6, V6uhu6, C7uhu6, J7uhu6, Q7uhu6, X7uhu6, E8uhu6, L8uhu6, S8uhu6, Z8uhu6;
wire G9uhu6, N9uhu6, U9uhu6, Bauhu6, Iauhu6, Pauhu6, Wauhu6, Dbuhu6, Kbuhu6, Rbuhu6;
wire Ybuhu6, Fcuhu6, Mcuhu6, Tcuhu6, Aduhu6, Hduhu6, Oduhu6, Vduhu6, Ceuhu6, Jeuhu6;
wire Qeuhu6, Xeuhu6, Efuhu6, Lfuhu6, Sfuhu6, Zfuhu6, Gguhu6, Nguhu6, Uguhu6, Bhuhu6;
wire Ihuhu6, Phuhu6, Whuhu6, Diuhu6, Kiuhu6, Riuhu6, Yiuhu6, Fjuhu6, Mjuhu6, Tjuhu6;
wire Akuhu6, Hkuhu6, Okuhu6, Vkuhu6, Cluhu6, Jluhu6, Qluhu6, Xluhu6, Emuhu6, Lmuhu6;
wire Smuhu6, Zmuhu6, Gnuhu6, Nnuhu6, Unuhu6, Bouhu6, Iouhu6, Pouhu6, Wouhu6, Dpuhu6;
wire Kpuhu6, Rpuhu6, Ypuhu6, Fquhu6, Mquhu6, Tquhu6, Aruhu6, Hruhu6, Oruhu6, Vruhu6;
wire Csuhu6, Jsuhu6, Qsuhu6, Xsuhu6, Etuhu6, Ltuhu6, Stuhu6, Ztuhu6, Guuhu6, Nuuhu6;
wire Uuuhu6, Bvuhu6, Ivuhu6, Pvuhu6, Wvuhu6, Dwuhu6, Kwuhu6, Rwuhu6, Ywuhu6, Fxuhu6;
wire Mxuhu6, Txuhu6, Ayuhu6, Hyuhu6, Oyuhu6, Vyuhu6, Czuhu6, Jzuhu6, Qzuhu6, Xzuhu6;
wire E0vhu6, L0vhu6, S0vhu6, Z0vhu6, G1vhu6, N1vhu6, U1vhu6, B2vhu6, I2vhu6, P2vhu6;
wire W2vhu6, D3vhu6, K3vhu6, R3vhu6, Y3vhu6, F4vhu6, M4vhu6, T4vhu6, A5vhu6, H5vhu6;
wire O5vhu6, V5vhu6, C6vhu6, J6vhu6, Q6vhu6, X6vhu6, E7vhu6, L7vhu6, S7vhu6, Z7vhu6;
wire G8vhu6, N8vhu6, U8vhu6, B9vhu6, I9vhu6, P9vhu6, W9vhu6, Davhu6, Kavhu6, Ravhu6;
wire Yavhu6, Fbvhu6, Mbvhu6, Tbvhu6, Acvhu6, Hcvhu6, Ocvhu6, Vcvhu6, Cdvhu6, Jdvhu6;
wire Qdvhu6, Xdvhu6, Eevhu6, Levhu6, Sevhu6, Zevhu6, Gfvhu6, Nfvhu6, Ufvhu6, Bgvhu6;
wire Igvhu6, Pgvhu6, Wgvhu6, Dhvhu6, Khvhu6, Rhvhu6, Yhvhu6, Fivhu6, Mivhu6, Tivhu6;
wire Ajvhu6, Hjvhu6, Ojvhu6, Vjvhu6, Ckvhu6, Jkvhu6, Qkvhu6, Xkvhu6, Elvhu6, Llvhu6;
wire Slvhu6, Zlvhu6, Gmvhu6, Nmvhu6, Umvhu6, Bnvhu6, Invhu6, Pnvhu6, Wnvhu6, Dovhu6;
wire Kovhu6, Rovhu6, Yovhu6, Fpvhu6, Mpvhu6, Tpvhu6, Aqvhu6, Hqvhu6, Oqvhu6, Vqvhu6;
wire Crvhu6, Jrvhu6, Qrvhu6, Xrvhu6, Esvhu6, Lsvhu6, Ssvhu6, Zsvhu6, Gtvhu6, Ntvhu6;
wire Utvhu6, Buvhu6, Iuvhu6, Puvhu6, Wuvhu6, Dvvhu6, Kvvhu6, Rvvhu6, Yvvhu6, Fwvhu6;
wire Mwvhu6, Twvhu6, Axvhu6, Hxvhu6, Oxvhu6, Vxvhu6, Cyvhu6, Jyvhu6, Qyvhu6, Xyvhu6;
wire Ezvhu6, Lzvhu6, Szvhu6, Zzvhu6, G0whu6, N0whu6, U0whu6, B1whu6, I1whu6, P1whu6;
wire W1whu6, D2whu6, K2whu6, R2whu6, Y2whu6, F3whu6, M3whu6, T3whu6, A4whu6, H4whu6;
wire O4whu6, V4whu6, C5whu6, J5whu6, Q5whu6, X5whu6, E6whu6, L6whu6, S6whu6, Z6whu6;
wire G7whu6, N7whu6, U7whu6, B8whu6, I8whu6, P8whu6, W8whu6, D9whu6, K9whu6, R9whu6;
wire Y9whu6, Fawhu6, Mawhu6, Tawhu6, Abwhu6, Hbwhu6, Obwhu6, Vbwhu6, Ccwhu6, Jcwhu6;
wire Qcwhu6, Xcwhu6, Edwhu6, Ldwhu6, Sdwhu6, Zdwhu6, Gewhu6, Newhu6, Uewhu6, Bfwhu6;
wire Ifwhu6, Pfwhu6, Wfwhu6, Dgwhu6, Kgwhu6, Rgwhu6, Ygwhu6, Fhwhu6, Mhwhu6, Thwhu6;
wire Aiwhu6, Hiwhu6, Oiwhu6, Viwhu6, Cjwhu6, Jjwhu6, Qjwhu6, Xjwhu6, Ekwhu6, Lkwhu6;
wire Skwhu6, Zkwhu6, Glwhu6, Nlwhu6, Ulwhu6, Bmwhu6, Imwhu6, Pmwhu6, Wmwhu6, Dnwhu6;
wire Knwhu6, Rnwhu6, Ynwhu6, Fowhu6, Mowhu6, Towhu6, Apwhu6, Hpwhu6, Opwhu6, Vpwhu6;
wire Cqwhu6, Jqwhu6, Qqwhu6, Xqwhu6, Erwhu6, Lrwhu6, Srwhu6, Zrwhu6, Gswhu6, Nswhu6;
wire Uswhu6, Btwhu6, Itwhu6, Ptwhu6, Wtwhu6, Duwhu6, Kuwhu6, Ruwhu6, Yuwhu6, Fvwhu6;
wire Mvwhu6, Tvwhu6, Awwhu6, Hwwhu6, Owwhu6, Vwwhu6, Cxwhu6, Jxwhu6, Qxwhu6, Xxwhu6;
wire Eywhu6, Lywhu6, Sywhu6, Zywhu6, Gzwhu6, Nzwhu6, Uzwhu6, B0xhu6, I0xhu6, P0xhu6;
wire W0xhu6, D1xhu6, K1xhu6, R1xhu6, Y1xhu6, F2xhu6, M2xhu6, T2xhu6, A3xhu6, H3xhu6;
wire O3xhu6, V3xhu6, C4xhu6, J4xhu6, Q4xhu6, X4xhu6, E5xhu6, L5xhu6, S5xhu6, Z5xhu6;
wire G6xhu6, N6xhu6, U6xhu6, B7xhu6, I7xhu6, P7xhu6, W7xhu6, D8xhu6, K8xhu6, R8xhu6;
wire Y8xhu6, F9xhu6, M9xhu6, T9xhu6, Aaxhu6, Haxhu6, Oaxhu6, Vaxhu6, Cbxhu6, Jbxhu6;
wire Qbxhu6, Xbxhu6, Ecxhu6, Lcxhu6, Scxhu6, Zcxhu6, Gdxhu6, Ndxhu6, Udxhu6, Bexhu6;
wire Iexhu6, Pexhu6, Wexhu6, Dfxhu6, Kfxhu6, Rfxhu6, Yfxhu6, Fgxhu6, Mgxhu6, Tgxhu6;
wire Ahxhu6, Hhxhu6, Ohxhu6, Vhxhu6, Cixhu6, Jixhu6, Qixhu6, Xixhu6, Ejxhu6, Ljxhu6;
wire Sjxhu6, Zjxhu6, Gkxhu6, Nkxhu6, Ukxhu6, Blxhu6, Ilxhu6, Plxhu6, Wlxhu6, Dmxhu6;
wire Kmxhu6, Rmxhu6, Ymxhu6, Fnxhu6, Mnxhu6, Tnxhu6, Aoxhu6, Hoxhu6, Ooxhu6, Voxhu6;
wire Cpxhu6, Jpxhu6, Qpxhu6, Xpxhu6, Eqxhu6, Lqxhu6, Sqxhu6, Zqxhu6, Grxhu6, Nrxhu6;
wire Urxhu6, Bsxhu6, Isxhu6, Psxhu6, Wsxhu6, Dtxhu6, Ktxhu6, Rtxhu6, Ytxhu6, Fuxhu6;
wire Muxhu6, Tuxhu6, Avxhu6, Hvxhu6, Ovxhu6, Vvxhu6, Cwxhu6, Jwxhu6, Qwxhu6, Xwxhu6;
wire Exxhu6, Lxxhu6, Sxxhu6, Zxxhu6, Gyxhu6, Nyxhu6, Uyxhu6, Bzxhu6, Izxhu6, Pzxhu6;
wire Wzxhu6, D0yhu6, K0yhu6, R0yhu6, Y0yhu6, F1yhu6, M1yhu6, T1yhu6, A2yhu6, H2yhu6;
wire O2yhu6, V2yhu6, C3yhu6, J3yhu6, Q3yhu6, X3yhu6, E4yhu6, L4yhu6, S4yhu6, Z4yhu6;
wire G5yhu6, N5yhu6, U5yhu6, B6yhu6, I6yhu6, P6yhu6, W6yhu6, D7yhu6, K7yhu6, R7yhu6;
wire Y7yhu6, F8yhu6, M8yhu6, T8yhu6, A9yhu6, H9yhu6, O9yhu6, V9yhu6, Cayhu6, Jayhu6;
wire Qayhu6, Xayhu6, Ebyhu6, Lbyhu6, Sbyhu6, Zbyhu6, Gcyhu6, Ncyhu6, Ucyhu6, Bdyhu6;
wire Idyhu6, Pdyhu6, Wdyhu6, Deyhu6, Keyhu6, Reyhu6, Yeyhu6, Ffyhu6, Mfyhu6, Tfyhu6;
wire Agyhu6, Hgyhu6, Ogyhu6, Vgyhu6, Chyhu6, Jhyhu6, Qhyhu6, Xhyhu6, Eiyhu6, Liyhu6;
wire Siyhu6, Ziyhu6, Gjyhu6, Njyhu6, Ujyhu6, Bkyhu6, Ikyhu6, Pkyhu6, Wkyhu6, Dlyhu6;
wire Klyhu6, Rlyhu6, Ylyhu6, Fmyhu6, Mmyhu6, Tmyhu6, Anyhu6, Hnyhu6, Onyhu6, Vnyhu6;
wire Coyhu6, Joyhu6, Qoyhu6, Xoyhu6, Epyhu6, Lpyhu6, Spyhu6, Zpyhu6, Gqyhu6, Nqyhu6;
wire Uqyhu6, Bryhu6, Iryhu6, Pryhu6, Wryhu6, Dsyhu6, Ksyhu6, Rsyhu6, Ysyhu6, Ftyhu6;
wire Mtyhu6, Ttyhu6, Auyhu6, Huyhu6, Ouyhu6, Vuyhu6, Cvyhu6, Jvyhu6, Qvyhu6, Xvyhu6;
wire Ewyhu6, Lwyhu6, Swyhu6, Zwyhu6, Gxyhu6, Nxyhu6, Uxyhu6, Byyhu6, Iyyhu6, Pyyhu6;
wire Wyyhu6, Dzyhu6, Kzyhu6, Rzyhu6, Yzyhu6, F0zhu6, M0zhu6, T0zhu6, A1zhu6, H1zhu6;
wire O1zhu6, V1zhu6, C2zhu6, J2zhu6, Q2zhu6, X2zhu6, E3zhu6, L3zhu6, S3zhu6, Z3zhu6;
wire G4zhu6, N4zhu6, U4zhu6, B5zhu6, I5zhu6, P5zhu6, W5zhu6, D6zhu6, K6zhu6, R6zhu6;
wire Y6zhu6, F7zhu6, M7zhu6, T7zhu6, A8zhu6, H8zhu6, O8zhu6, V8zhu6, C9zhu6, J9zhu6;
wire Q9zhu6, X9zhu6, Eazhu6, Lazhu6, Sazhu6, Zazhu6, Gbzhu6, Nbzhu6, Ubzhu6, Bczhu6;
wire Iczhu6, Pczhu6, Wczhu6, Ddzhu6, Kdzhu6, Rdzhu6, Ydzhu6, Fezhu6, Mezhu6, Tezhu6;
wire Afzhu6, Hfzhu6, Ofzhu6, Vfzhu6, Cgzhu6, Jgzhu6, Qgzhu6, Xgzhu6, Ehzhu6, Lhzhu6;
wire Shzhu6, Zhzhu6, Gizhu6, Nizhu6, Uizhu6, Bjzhu6, Ijzhu6, Pjzhu6, Wjzhu6, Dkzhu6;
wire Kkzhu6, Rkzhu6, Ykzhu6, Flzhu6, Mlzhu6, Tlzhu6, Amzhu6, Hmzhu6, Omzhu6, Vmzhu6;
wire Cnzhu6, Jnzhu6, Qnzhu6, Xnzhu6, Eozhu6, Lozhu6, Sozhu6, Zozhu6, Gpzhu6, Npzhu6;
wire Upzhu6, Bqzhu6, Iqzhu6, Pqzhu6, Wqzhu6, Drzhu6, Krzhu6, Rrzhu6, Yrzhu6, Fszhu6;
wire Mszhu6, Tszhu6, Atzhu6, Htzhu6, Otzhu6, Vtzhu6, Cuzhu6, Juzhu6, Quzhu6, Xuzhu6;
wire Evzhu6, Lvzhu6, Svzhu6, Zvzhu6, Gwzhu6, Nwzhu6, Uwzhu6, Bxzhu6, Ixzhu6, Pxzhu6;
wire Wxzhu6, Dyzhu6, Kyzhu6, Ryzhu6, Yyzhu6, Fzzhu6, Mzzhu6, Tzzhu6, A00iu6, H00iu6;
wire O00iu6, V00iu6, C10iu6, J10iu6, Q10iu6, X10iu6, E20iu6, L20iu6, S20iu6, Z20iu6;
wire G30iu6, N30iu6, U30iu6, B40iu6, I40iu6, P40iu6, W40iu6, D50iu6, K50iu6, R50iu6;
wire Y50iu6, F60iu6, M60iu6, T60iu6, A70iu6, H70iu6, O70iu6, V70iu6, C80iu6, J80iu6;
wire Q80iu6, X80iu6, E90iu6, L90iu6, S90iu6, Z90iu6, Ga0iu6, Na0iu6, Ua0iu6, Bb0iu6;
wire Ib0iu6, Pb0iu6, Wb0iu6, Dc0iu6, Kc0iu6, Rc0iu6, Yc0iu6, Fd0iu6, Md0iu6, Td0iu6;
wire Ae0iu6, He0iu6, Oe0iu6, Ve0iu6, Cf0iu6, Jf0iu6, Qf0iu6, Xf0iu6, Eg0iu6, Lg0iu6;
wire Sg0iu6, Zg0iu6, Gh0iu6, Nh0iu6, Uh0iu6, Bi0iu6, Ii0iu6, Pi0iu6, Wi0iu6, Dj0iu6;
wire Kj0iu6, Rj0iu6, Yj0iu6, Fk0iu6, Mk0iu6, Tk0iu6, Al0iu6, Hl0iu6, Ol0iu6, Vl0iu6;
wire Cm0iu6, Jm0iu6, Qm0iu6, Xm0iu6, En0iu6, Ln0iu6, Sn0iu6, Zn0iu6, Go0iu6, No0iu6;
wire Uo0iu6, Bp0iu6, Ip0iu6, Pp0iu6, Wp0iu6, Dq0iu6, Kq0iu6, Rq0iu6, Yq0iu6, Fr0iu6;
wire Mr0iu6, Tr0iu6, As0iu6, Hs0iu6, Os0iu6, Vs0iu6, Ct0iu6, Jt0iu6, Qt0iu6, Xt0iu6;
wire Eu0iu6, Lu0iu6, Su0iu6, Zu0iu6, Gv0iu6, Nv0iu6, Uv0iu6, Bw0iu6, Iw0iu6, Pw0iu6;
wire Ww0iu6, Dx0iu6, Kx0iu6, Rx0iu6, Yx0iu6, Fy0iu6, My0iu6, Ty0iu6, Az0iu6, Hz0iu6;
wire Oz0iu6, Vz0iu6, C01iu6, J01iu6, Q01iu6, X01iu6, E11iu6, L11iu6, S11iu6, Z11iu6;
wire G21iu6, N21iu6, U21iu6, B31iu6, I31iu6, P31iu6, W31iu6, D41iu6, K41iu6, R41iu6;
wire Y41iu6, F51iu6, M51iu6, T51iu6, A61iu6, H61iu6, O61iu6, V61iu6, C71iu6, J71iu6;
wire Q71iu6, X71iu6, E81iu6, L81iu6, S81iu6, Z81iu6, G91iu6, N91iu6, U91iu6, Ba1iu6;
wire Ia1iu6, Pa1iu6, Wa1iu6, Db1iu6, Kb1iu6, Rb1iu6, Yb1iu6, Fc1iu6, Mc1iu6, Tc1iu6;
wire Ad1iu6, Hd1iu6, Od1iu6, Vd1iu6, Ce1iu6, Je1iu6, Qe1iu6, Xe1iu6, Ef1iu6, Lf1iu6;
wire Sf1iu6, Zf1iu6, Gg1iu6, Ng1iu6, Ug1iu6, Bh1iu6, Ih1iu6, Ph1iu6, Wh1iu6, Di1iu6;
wire Ki1iu6, Ri1iu6, Yi1iu6, Fj1iu6, Mj1iu6, Tj1iu6, Ak1iu6, Hk1iu6, Ok1iu6, Vk1iu6;
wire Cl1iu6, Jl1iu6, Ql1iu6, Xl1iu6, Em1iu6, Lm1iu6, Sm1iu6, Zm1iu6, Gn1iu6, Nn1iu6;
wire Un1iu6, Bo1iu6, Io1iu6, Po1iu6, Wo1iu6, Dp1iu6, Kp1iu6, Rp1iu6, Yp1iu6, Fq1iu6;
wire Mq1iu6, Tq1iu6, Ar1iu6, Hr1iu6, Or1iu6, Vr1iu6, Cs1iu6, Js1iu6, Qs1iu6, Xs1iu6;
wire Et1iu6, Lt1iu6, St1iu6, Zt1iu6, Gu1iu6, Nu1iu6, Uu1iu6, Bv1iu6, Iv1iu6, Pv1iu6;
wire Wv1iu6, Dw1iu6, Kw1iu6, Rw1iu6, Yw1iu6, Fx1iu6, Mx1iu6, Tx1iu6, Ay1iu6, Hy1iu6;
wire Oy1iu6, Vy1iu6, Cz1iu6, Jz1iu6, Qz1iu6, Xz1iu6, E02iu6, L02iu6, S02iu6, Z02iu6;
wire G12iu6, N12iu6, U12iu6, B22iu6, I22iu6, P22iu6, W22iu6, D32iu6, K32iu6, R32iu6;
wire Y32iu6, F42iu6, M42iu6, T42iu6, A52iu6, H52iu6, O52iu6, V52iu6, C62iu6, J62iu6;
wire Q62iu6, X62iu6, E72iu6, L72iu6, S72iu6, Z72iu6, G82iu6, N82iu6, U82iu6, B92iu6;
wire I92iu6, P92iu6, W92iu6, Da2iu6, Ka2iu6, Ra2iu6, Ya2iu6, Fb2iu6, Mb2iu6, Tb2iu6;
wire Ac2iu6, Hc2iu6, Oc2iu6, Vc2iu6, Cd2iu6, Jd2iu6, Qd2iu6, Xd2iu6, Ee2iu6, Le2iu6;
wire Se2iu6, Ze2iu6, Gf2iu6, Nf2iu6, Uf2iu6, Bg2iu6, Ig2iu6, Pg2iu6, Wg2iu6, Dh2iu6;
wire Kh2iu6, Rh2iu6, Yh2iu6, Fi2iu6, Mi2iu6, Ti2iu6, Aj2iu6, Hj2iu6, Oj2iu6, Vj2iu6;
wire Ck2iu6, Jk2iu6, Qk2iu6, Xk2iu6, El2iu6, Ll2iu6, Sl2iu6, Zl2iu6, Gm2iu6, Nm2iu6;
wire Um2iu6, Bn2iu6, In2iu6, Pn2iu6, Wn2iu6, Do2iu6, Ko2iu6, Ro2iu6, Yo2iu6, Fp2iu6;
wire Mp2iu6, Tp2iu6, Aq2iu6, Hq2iu6, Oq2iu6, Vq2iu6, Cr2iu6, Jr2iu6, Qr2iu6, Xr2iu6;
wire Es2iu6, Ls2iu6, Ss2iu6, Zs2iu6, Gt2iu6, Nt2iu6, Ut2iu6, Bu2iu6, Iu2iu6, Pu2iu6;
wire Wu2iu6, Dv2iu6, Kv2iu6, Rv2iu6, Yv2iu6, Fw2iu6, Mw2iu6, Tw2iu6, Ax2iu6, Hx2iu6;
wire Ox2iu6, Vx2iu6, Cy2iu6, Jy2iu6, Qy2iu6, Xy2iu6, Ez2iu6, Lz2iu6, Sz2iu6, Zz2iu6;
wire G03iu6, N03iu6, U03iu6, B13iu6, I13iu6, P13iu6, W13iu6, D23iu6, K23iu6, R23iu6;
wire Y23iu6, F33iu6, M33iu6, T33iu6, A43iu6, H43iu6, O43iu6, V43iu6, C53iu6, J53iu6;
wire Q53iu6, X53iu6, E63iu6, L63iu6, S63iu6, Z63iu6, G73iu6, N73iu6, U73iu6, B83iu6;
wire I83iu6, P83iu6, W83iu6, D93iu6, K93iu6, R93iu6, Y93iu6, Fa3iu6, Ma3iu6, Ta3iu6;
wire Ab3iu6, Hb3iu6, Ob3iu6, Vb3iu6, Cc3iu6, Jc3iu6, Qc3iu6, Xc3iu6, Ed3iu6, Ld3iu6;
wire Sd3iu6, Zd3iu6, Ge3iu6, Ne3iu6, Ue3iu6, Bf3iu6, If3iu6, Pf3iu6, Wf3iu6, Dg3iu6;
wire Kg3iu6, Rg3iu6, Yg3iu6, Fh3iu6, Mh3iu6, Th3iu6, Ai3iu6, Hi3iu6, Oi3iu6, Vi3iu6;
wire Cj3iu6, Jj3iu6, Qj3iu6, Xj3iu6, Ek3iu6, Lk3iu6, Sk3iu6, Zk3iu6, Gl3iu6, Nl3iu6;
wire Ul3iu6, Bm3iu6, Im3iu6, Pm3iu6, Wm3iu6, Dn3iu6, Kn3iu6, Rn3iu6, Yn3iu6, Fo3iu6;
wire Mo3iu6, To3iu6, Ap3iu6, Hp3iu6, Op3iu6, Vp3iu6, Cq3iu6, Jq3iu6, Qq3iu6, Xq3iu6;
wire Er3iu6, Lr3iu6, Sr3iu6, Zr3iu6, Gs3iu6, Ns3iu6, Us3iu6, Bt3iu6, It3iu6, Pt3iu6;
wire Wt3iu6, Du3iu6, Ku3iu6, Ru3iu6, Yu3iu6, Fv3iu6, Mv3iu6, Tv3iu6, Aw3iu6, Hw3iu6;
wire Ow3iu6, Vw3iu6, Cx3iu6, Jx3iu6, Qx3iu6, Xx3iu6, Ey3iu6, Ly3iu6, Sy3iu6, Zy3iu6;
wire Gz3iu6, Nz3iu6, Uz3iu6, B04iu6, I04iu6, P04iu6, W04iu6, D14iu6, K14iu6, R14iu6;
wire Y14iu6, F24iu6, M24iu6, T24iu6, A34iu6, H34iu6, O34iu6, V34iu6, C44iu6, J44iu6;
wire Q44iu6, X44iu6, E54iu6, L54iu6, S54iu6, Z54iu6, G64iu6, N64iu6, U64iu6, B74iu6;
wire I74iu6, P74iu6, W74iu6, D84iu6, K84iu6, R84iu6, Y84iu6, F94iu6, M94iu6, T94iu6;
wire Aa4iu6, Ha4iu6, Oa4iu6, Va4iu6, Cb4iu6, Jb4iu6, Qb4iu6, Xb4iu6, Ec4iu6, Lc4iu6;
wire Sc4iu6, Zc4iu6, Gd4iu6, Nd4iu6, Ud4iu6, Be4iu6, Ie4iu6, Pe4iu6, We4iu6, Df4iu6;
wire Kf4iu6, Rf4iu6, Yf4iu6, Fg4iu6, Mg4iu6, Tg4iu6, Ah4iu6, Hh4iu6, Oh4iu6, Vh4iu6;
wire Ci4iu6, Ji4iu6, Qi4iu6, Xi4iu6, Ej4iu6, Lj4iu6, Sj4iu6, Zj4iu6, Gk4iu6, Nk4iu6;
wire Uk4iu6, Bl4iu6, Il4iu6, Pl4iu6, Wl4iu6, Dm4iu6, Km4iu6, Rm4iu6, Ym4iu6, Fn4iu6;
wire Mn4iu6, Tn4iu6, Ao4iu6, Ho4iu6, Oo4iu6, Vo4iu6, Cp4iu6, Jp4iu6, Qp4iu6, Xp4iu6;
wire Eq4iu6, Lq4iu6, Sq4iu6, Zq4iu6, Gr4iu6, Nr4iu6, Ur4iu6, Bs4iu6, Is4iu6, Ps4iu6;
wire Ws4iu6, Dt4iu6, Kt4iu6, Rt4iu6, Yt4iu6, Fu4iu6, Mu4iu6, Tu4iu6, Av4iu6, Hv4iu6;
wire Ov4iu6, Vv4iu6, Cw4iu6, Jw4iu6, Qw4iu6, Xw4iu6, Ex4iu6, Lx4iu6, Sx4iu6, Zx4iu6;
wire Gy4iu6, Ny4iu6, Uy4iu6, Bz4iu6, Iz4iu6, Pz4iu6, Wz4iu6, D05iu6, K05iu6, R05iu6;
wire Y05iu6, F15iu6, M15iu6, T15iu6, A25iu6, H25iu6, O25iu6, V25iu6, C35iu6, J35iu6;
wire Q35iu6, X35iu6, E45iu6, L45iu6, S45iu6, Z45iu6, G55iu6, N55iu6, U55iu6, B65iu6;
wire I65iu6, P65iu6, W65iu6, D75iu6, K75iu6, R75iu6, Y75iu6, F85iu6, M85iu6, T85iu6;
wire A95iu6, H95iu6, O95iu6, V95iu6, Ca5iu6, Ja5iu6, Qa5iu6, Xa5iu6, Eb5iu6, Lb5iu6;
wire Sb5iu6, Zb5iu6, Gc5iu6, Nc5iu6, Uc5iu6, Bd5iu6, Id5iu6, Pd5iu6, Wd5iu6, De5iu6;
wire Ke5iu6, Re5iu6, Ye5iu6, Ff5iu6, Mf5iu6, Tf5iu6, Ag5iu6, Hg5iu6, Og5iu6, Vg5iu6;
wire Ch5iu6, Jh5iu6, Qh5iu6, Xh5iu6, Ei5iu6, Li5iu6, Si5iu6, Zi5iu6, Gj5iu6, Nj5iu6;
wire Uj5iu6, Bk5iu6, Ik5iu6, Pk5iu6, Wk5iu6, Dl5iu6, Kl5iu6, Rl5iu6, Yl5iu6, Fm5iu6;
wire Mm5iu6, Tm5iu6, An5iu6, Hn5iu6, On5iu6, Vn5iu6, Co5iu6, Jo5iu6, Qo5iu6, Xo5iu6;
wire Ep5iu6, Lp5iu6, Sp5iu6, Zp5iu6, Gq5iu6, Nq5iu6, Uq5iu6, Br5iu6, Ir5iu6, Pr5iu6;
wire Wr5iu6, Ds5iu6, Ks5iu6, Rs5iu6, Ys5iu6, Ft5iu6, Mt5iu6, Tt5iu6, Au5iu6, Hu5iu6;
wire Ou5iu6, Vu5iu6, Cv5iu6, Jv5iu6, Qv5iu6, Xv5iu6, Ew5iu6, Lw5iu6, Sw5iu6, Zw5iu6;
wire Gx5iu6, Nx5iu6, Ux5iu6, By5iu6, Iy5iu6, Py5iu6, Wy5iu6, Dz5iu6, Kz5iu6, Rz5iu6;
wire Yz5iu6, F06iu6, M06iu6, T06iu6, A16iu6, H16iu6, O16iu6, V16iu6, C26iu6, J26iu6;
wire Q26iu6, X26iu6, E36iu6, L36iu6, S36iu6, Z36iu6, G46iu6, N46iu6, U46iu6, B56iu6;
wire I56iu6, P56iu6, W56iu6, D66iu6, K66iu6, R66iu6, Y66iu6, F76iu6, M76iu6, T76iu6;
wire A86iu6, H86iu6, O86iu6, V86iu6, C96iu6, J96iu6, Q96iu6, X96iu6, Ea6iu6, La6iu6;
wire Sa6iu6, Za6iu6, Gb6iu6, Nb6iu6, Ub6iu6, Bc6iu6, Ic6iu6, Pc6iu6, Wc6iu6, Dd6iu6;
wire Kd6iu6, Rd6iu6, Yd6iu6, Fe6iu6, Me6iu6, Te6iu6, Af6iu6, Hf6iu6, Of6iu6, Vf6iu6;
wire Cg6iu6, Jg6iu6, Qg6iu6, Xg6iu6, Eh6iu6, Lh6iu6, Sh6iu6, Zh6iu6, Gi6iu6, Ni6iu6;
wire Ui6iu6, Bj6iu6, Ij6iu6, Pj6iu6, Wj6iu6, Dk6iu6, Kk6iu6, Rk6iu6, Yk6iu6, Fl6iu6;
wire Ml6iu6, Tl6iu6, Am6iu6, Hm6iu6, Om6iu6, Vm6iu6, Cn6iu6, Jn6iu6, Qn6iu6, Xn6iu6;
wire Eo6iu6, Lo6iu6, So6iu6, Zo6iu6, Gp6iu6, Np6iu6, Up6iu6, Bq6iu6, Iq6iu6, Pq6iu6;
wire Wq6iu6, Dr6iu6, Kr6iu6, Rr6iu6, Yr6iu6, Fs6iu6, Ms6iu6, Ts6iu6, At6iu6, Ht6iu6;
wire Ot6iu6, Vt6iu6, Cu6iu6, Ju6iu6, Qu6iu6, Xu6iu6, Ev6iu6, Lv6iu6, Sv6iu6, Zv6iu6;
wire Gw6iu6, Nw6iu6, Uw6iu6, Bx6iu6, Ix6iu6, Px6iu6, Wx6iu6, Dy6iu6, Ky6iu6, Ry6iu6;
wire Yy6iu6, Fz6iu6, Mz6iu6, Tz6iu6, A07iu6, H07iu6, O07iu6, V07iu6, C17iu6, J17iu6;
wire Q17iu6, X17iu6, E27iu6, L27iu6, S27iu6, Z27iu6, G37iu6, N37iu6, U37iu6, B47iu6;
wire I47iu6, P47iu6, W47iu6, D57iu6, K57iu6, R57iu6, Y57iu6, F67iu6, M67iu6, T67iu6;
wire A77iu6, H77iu6, O77iu6, V77iu6, C87iu6, J87iu6, Q87iu6, X87iu6, E97iu6, L97iu6;
wire S97iu6, Z97iu6, Ga7iu6, Na7iu6, Ua7iu6, Bb7iu6, Ib7iu6, Pb7iu6, Wb7iu6, Dc7iu6;
wire Kc7iu6, Rc7iu6, Yc7iu6, Fd7iu6, Md7iu6, Td7iu6, Ae7iu6, He7iu6, Oe7iu6, Ve7iu6;
wire Cf7iu6, Jf7iu6, Qf7iu6, Xf7iu6, Eg7iu6, Lg7iu6, Sg7iu6, Zg7iu6, Gh7iu6, Nh7iu6;
wire Uh7iu6, Bi7iu6, Ii7iu6, Pi7iu6, Wi7iu6, Dj7iu6, Kj7iu6, Rj7iu6, Yj7iu6, Fk7iu6;
wire Mk7iu6, Tk7iu6, Al7iu6, Hl7iu6, Ol7iu6, Vl7iu6, Cm7iu6, Jm7iu6, Qm7iu6, Xm7iu6;
wire En7iu6, Ln7iu6, Sn7iu6, Zn7iu6, Go7iu6, No7iu6, Uo7iu6, Bp7iu6, Ip7iu6, Pp7iu6;
wire Wp7iu6, Dq7iu6, Kq7iu6, Rq7iu6, Yq7iu6, Fr7iu6, Mr7iu6, Tr7iu6, As7iu6, Hs7iu6;
wire Os7iu6, Vs7iu6, Ct7iu6, Jt7iu6, Qt7iu6, Xt7iu6, Eu7iu6, Lu7iu6, Su7iu6, Zu7iu6;
wire Gv7iu6, Nv7iu6, Uv7iu6, Bw7iu6, Iw7iu6, Pw7iu6, Ww7iu6, Dx7iu6, Kx7iu6, Rx7iu6;
wire Yx7iu6, Fy7iu6, My7iu6, Ty7iu6, Az7iu6, Hz7iu6, Oz7iu6, Vz7iu6, C08iu6, J08iu6;
wire Q08iu6, X08iu6, E18iu6, L18iu6, S18iu6, Z18iu6, G28iu6, N28iu6, U28iu6, B38iu6;
wire I38iu6, P38iu6, W38iu6, D48iu6, K48iu6, R48iu6, Y48iu6, F58iu6, M58iu6, T58iu6;
wire A68iu6, H68iu6, O68iu6, V68iu6, C78iu6, J78iu6, Q78iu6, X78iu6, E88iu6, L88iu6;
wire S88iu6, Z88iu6, G98iu6, N98iu6, U98iu6, Ba8iu6, Ia8iu6, Pa8iu6, Wa8iu6, Db8iu6;
wire Kb8iu6, Rb8iu6, Yb8iu6, Fc8iu6, Mc8iu6, Tc8iu6, Ad8iu6, Hd8iu6, Od8iu6, Vd8iu6;
wire Ce8iu6, Je8iu6, Qe8iu6, Xe8iu6, Ef8iu6, Lf8iu6, Sf8iu6, Zf8iu6, Gg8iu6, Ng8iu6;
wire Ug8iu6, Bh8iu6, Ih8iu6, Ph8iu6, Wh8iu6, Di8iu6, Ki8iu6, Ri8iu6, Yi8iu6, Fj8iu6;
wire Mj8iu6, Tj8iu6, Ak8iu6, Hk8iu6, Ok8iu6, Vk8iu6, Cl8iu6, Jl8iu6, Ql8iu6, Xl8iu6;
wire Em8iu6, Lm8iu6, Sm8iu6, Zm8iu6, Gn8iu6, Nn8iu6, Un8iu6, Bo8iu6, Io8iu6, Po8iu6;
wire Wo8iu6, Dp8iu6, Kp8iu6, Rp8iu6, Yp8iu6, Fq8iu6, Mq8iu6, Tq8iu6, Ar8iu6, Hr8iu6;
wire Or8iu6, Vr8iu6, Cs8iu6, Js8iu6, Qs8iu6, Xs8iu6, Et8iu6, Lt8iu6, St8iu6, Zt8iu6;
wire Gu8iu6, Nu8iu6, Uu8iu6, Bv8iu6, Iv8iu6, Pv8iu6, Wv8iu6, Dw8iu6, Kw8iu6, Rw8iu6;
wire Yw8iu6, Fx8iu6, Mx8iu6, Tx8iu6, Ay8iu6, Hy8iu6, Oy8iu6, Vy8iu6, Cz8iu6, Jz8iu6;
wire Qz8iu6, Xz8iu6, E09iu6, L09iu6, S09iu6, Z09iu6, G19iu6, N19iu6, U19iu6, B29iu6;
wire I29iu6, P29iu6, W29iu6, D39iu6, K39iu6, R39iu6, Y39iu6, F49iu6, M49iu6, T49iu6;
wire A59iu6, H59iu6, O59iu6, V59iu6, C69iu6, J69iu6, Q69iu6, X69iu6, E79iu6, L79iu6;
wire S79iu6, Z79iu6, G89iu6, N89iu6, U89iu6, B99iu6, I99iu6, P99iu6, W99iu6, Da9iu6;
wire Ka9iu6, Ra9iu6, Ya9iu6, Fb9iu6, Mb9iu6, Tb9iu6, Ac9iu6, Hc9iu6, Oc9iu6, Vc9iu6;
wire Cd9iu6, Jd9iu6, Qd9iu6, Xd9iu6, Ee9iu6, Le9iu6, Se9iu6, Ze9iu6, Gf9iu6, Nf9iu6;
wire Uf9iu6, Bg9iu6, Ig9iu6, Pg9iu6, Wg9iu6, Dh9iu6, Kh9iu6, Rh9iu6, Yh9iu6, Fi9iu6;
wire Mi9iu6, Ti9iu6, Aj9iu6, Hj9iu6, Oj9iu6, Vj9iu6, Ck9iu6, Jk9iu6, Qk9iu6, Xk9iu6;
wire El9iu6, Ll9iu6, Sl9iu6, Zl9iu6, Gm9iu6, Nm9iu6, Um9iu6, Bn9iu6, In9iu6, Pn9iu6;
wire Wn9iu6, Do9iu6, Ko9iu6, Ro9iu6, Yo9iu6, Fp9iu6, Mp9iu6, Tp9iu6, Aq9iu6, Hq9iu6;
wire Oq9iu6, Vq9iu6, Cr9iu6, Jr9iu6, Qr9iu6, Xr9iu6, Es9iu6, Ls9iu6, Ss9iu6, Zs9iu6;
wire Gt9iu6, Nt9iu6, Ut9iu6, Bu9iu6, Iu9iu6, Pu9iu6, Wu9iu6, Dv9iu6, Kv9iu6, Rv9iu6;
wire Yv9iu6, Fw9iu6, Mw9iu6, Tw9iu6, Ax9iu6, Hx9iu6, Ox9iu6, Vx9iu6, Cy9iu6, Jy9iu6;
wire Qy9iu6, Xy9iu6, Ez9iu6, Lz9iu6, Sz9iu6, Zz9iu6, G0aiu6, N0aiu6, U0aiu6, B1aiu6;
wire I1aiu6, P1aiu6, W1aiu6, D2aiu6, K2aiu6, R2aiu6, Y2aiu6, F3aiu6, M3aiu6, T3aiu6;
wire A4aiu6, H4aiu6, O4aiu6, V4aiu6, C5aiu6, J5aiu6, Q5aiu6, X5aiu6, E6aiu6, L6aiu6;
wire S6aiu6, Z6aiu6, G7aiu6, N7aiu6, U7aiu6, B8aiu6, I8aiu6, P8aiu6, W8aiu6, D9aiu6;
wire K9aiu6, R9aiu6, Y9aiu6, Faaiu6, Maaiu6, Taaiu6, Abaiu6, Hbaiu6, Obaiu6, Vbaiu6;
wire Ccaiu6, Jcaiu6, Qcaiu6, Xcaiu6, Edaiu6, Ldaiu6, Sdaiu6, Zdaiu6, Geaiu6, Neaiu6;
wire Ueaiu6, Bfaiu6, Ifaiu6, Pfaiu6, Wfaiu6, Dgaiu6, Kgaiu6, Rgaiu6, Ygaiu6, Fhaiu6;
wire Mhaiu6, Thaiu6, Aiaiu6, Hiaiu6, Oiaiu6, Viaiu6, Cjaiu6, Jjaiu6, Qjaiu6, Xjaiu6;
wire Ekaiu6, Lkaiu6, Skaiu6, Zkaiu6, Glaiu6, Nlaiu6, Ulaiu6, Bmaiu6, Imaiu6, Pmaiu6;
wire Wmaiu6, Dnaiu6, Knaiu6, Rnaiu6, Ynaiu6, Foaiu6, Moaiu6, Toaiu6, Apaiu6, Hpaiu6;
wire Opaiu6, Vpaiu6, Cqaiu6, Jqaiu6, Qqaiu6, Xqaiu6, Eraiu6, Lraiu6, Sraiu6, Zraiu6;
wire Gsaiu6, Nsaiu6, Usaiu6, Btaiu6, Itaiu6, Ptaiu6, Wtaiu6, Duaiu6, Kuaiu6, Ruaiu6;
wire Yuaiu6, Fvaiu6, Mvaiu6, Tvaiu6, Awaiu6, Hwaiu6, Owaiu6, Vwaiu6, Cxaiu6, Jxaiu6;
wire Qxaiu6, Xxaiu6, Eyaiu6, Lyaiu6, Syaiu6, Zyaiu6, Gzaiu6, Nzaiu6, Uzaiu6, B0biu6;
wire I0biu6, P0biu6, W0biu6, D1biu6, K1biu6, R1biu6, Y1biu6, F2biu6, M2biu6, T2biu6;
wire A3biu6, H3biu6, O3biu6, V3biu6, C4biu6, J4biu6, Q4biu6, X4biu6, E5biu6, L5biu6;
wire S5biu6, Z5biu6, G6biu6, N6biu6, U6biu6, B7biu6, I7biu6, P7biu6, W7biu6, D8biu6;
wire K8biu6, R8biu6, Y8biu6, F9biu6, M9biu6, T9biu6, Aabiu6, Habiu6, Oabiu6, Vabiu6;
wire Cbbiu6, Jbbiu6, Qbbiu6, Xbbiu6, Ecbiu6, Lcbiu6, Scbiu6, Zcbiu6, Gdbiu6, Ndbiu6;
wire Udbiu6, Bebiu6, Iebiu6, Pebiu6, Webiu6, Dfbiu6, Kfbiu6, Rfbiu6, Yfbiu6, Fgbiu6;
wire Mgbiu6, Tgbiu6, Ahbiu6, Hhbiu6, Ohbiu6, Vhbiu6, Cibiu6, Jibiu6, Qibiu6, Xibiu6;
wire Ejbiu6, Ljbiu6, Sjbiu6, Zjbiu6, Gkbiu6, Nkbiu6, Ukbiu6, Blbiu6, Ilbiu6, Plbiu6;
wire Wlbiu6, Dmbiu6, Kmbiu6, Rmbiu6, Ymbiu6, Fnbiu6, Mnbiu6, Tnbiu6, Aobiu6, Hobiu6;
wire Oobiu6, Vobiu6, Cpbiu6, Jpbiu6, Qpbiu6, Xpbiu6, Eqbiu6, Lqbiu6, Sqbiu6, Zqbiu6;
wire Grbiu6, Nrbiu6, Urbiu6, Bsbiu6, Isbiu6, Psbiu6, Wsbiu6, Dtbiu6, Ktbiu6, Rtbiu6;
wire Ytbiu6, Fubiu6, Mubiu6, Tubiu6, Avbiu6, Hvbiu6, Ovbiu6, Vvbiu6, Cwbiu6, Jwbiu6;
wire Qwbiu6, Xwbiu6, Exbiu6, Lxbiu6, Sxbiu6, Zxbiu6, Gybiu6, Nybiu6, Uybiu6, Bzbiu6;
wire Izbiu6, Pzbiu6, Wzbiu6, D0ciu6, K0ciu6, R0ciu6, Y0ciu6, F1ciu6, M1ciu6, T1ciu6;
wire A2ciu6, H2ciu6, O2ciu6, V2ciu6, C3ciu6, J3ciu6, Q3ciu6, X3ciu6, E4ciu6, L4ciu6;
wire S4ciu6, Z4ciu6, G5ciu6, N5ciu6, U5ciu6, B6ciu6, I6ciu6, P6ciu6, W6ciu6, D7ciu6;
wire K7ciu6, R7ciu6, Y7ciu6, F8ciu6, M8ciu6, T8ciu6, A9ciu6, H9ciu6, O9ciu6, V9ciu6;
wire Caciu6, Jaciu6, Qaciu6, Xaciu6, Ebciu6, Lbciu6, Sbciu6, Zbciu6, Gcciu6, Ncciu6;
wire Ucciu6, Bdciu6, Idciu6, Pdciu6, Wdciu6, Deciu6, Keciu6, Reciu6, Yeciu6, Ffciu6;
wire Mfciu6, Tfciu6, Agciu6, Hgciu6, Ogciu6, Vgciu6, Chciu6, Jhciu6, Qhciu6, Xhciu6;
wire Eiciu6, Liciu6, Siciu6, Ziciu6, Gjciu6, Njciu6, Ujciu6, Bkciu6, Ikciu6, Pkciu6;
wire Wkciu6, Dlciu6, Klciu6, Rlciu6, Ylciu6, Fmciu6, Mmciu6, Tmciu6, Anciu6, Hnciu6;
wire Onciu6, Vnciu6, Cociu6, Jociu6, Qociu6, Xociu6, Epciu6, Lpciu6, Spciu6, Zpciu6;
wire Gqciu6, Nqciu6, Uqciu6, Brciu6, Irciu6, Prciu6, Wrciu6, Dsciu6, Ksciu6, Rsciu6;
wire Ysciu6, Ftciu6, Mtciu6, Ttciu6, Auciu6, Huciu6, Ouciu6, Vuciu6, Cvciu6, Jvciu6;
wire Qvciu6, Xvciu6, Ewciu6, Lwciu6, Swciu6, Zwciu6, Gxciu6, Nxciu6, Uxciu6, Byciu6;
wire Iyciu6, Pyciu6, Wyciu6, Dzciu6, Kzciu6, Rzciu6, Yzciu6, F0diu6, M0diu6, T0diu6;
wire A1diu6, H1diu6, O1diu6, V1diu6, C2diu6, J2diu6, Q2diu6, X2diu6, E3diu6, L3diu6;
wire S3diu6, Z3diu6, G4diu6, N4diu6, U4diu6, B5diu6, I5diu6, P5diu6, W5diu6, D6diu6;
wire K6diu6, R6diu6, Y6diu6, F7diu6, M7diu6, T7diu6, A8diu6, H8diu6, O8diu6, V8diu6;
wire C9diu6, J9diu6, Q9diu6, X9diu6, Eadiu6, Ladiu6, Sadiu6, Zadiu6, Gbdiu6, Nbdiu6;
wire Ubdiu6, Bcdiu6, Icdiu6, Pcdiu6, Wcdiu6, Dddiu6, Kddiu6, Rddiu6, Yddiu6, Fediu6;
wire Mediu6, Tediu6, Afdiu6, Hfdiu6, Ofdiu6, Vfdiu6, Cgdiu6, Jgdiu6, Qgdiu6, Xgdiu6;
wire Ehdiu6, Lhdiu6, Shdiu6, Zhdiu6, Gidiu6, Nidiu6, Uidiu6, Bjdiu6, Ijdiu6, Pjdiu6;
wire Wjdiu6, Dkdiu6, Kkdiu6, Rkdiu6, Ykdiu6, Fldiu6, Mldiu6, Tldiu6, Amdiu6, Hmdiu6;
wire Omdiu6, Vmdiu6, Cndiu6, Jndiu6, Qndiu6, Xndiu6, Eodiu6, Lodiu6, Sodiu6, Zodiu6;
wire Gpdiu6, Npdiu6, Updiu6, Bqdiu6, Iqdiu6, Pqdiu6, Wqdiu6, Drdiu6, Krdiu6, Rrdiu6;
wire Yrdiu6, Fsdiu6, Msdiu6, Tsdiu6, Atdiu6, Htdiu6, Otdiu6, Vtdiu6, Cudiu6, Judiu6;
wire Qudiu6, Xudiu6, Evdiu6, Lvdiu6, Svdiu6, Zvdiu6, Gwdiu6, Nwdiu6, Uwdiu6, Bxdiu6;
wire Ixdiu6, Pxdiu6, Wxdiu6, Dydiu6, Kydiu6, Rydiu6, Yydiu6, Fzdiu6, Mzdiu6, Tzdiu6;
wire A0eiu6, H0eiu6, O0eiu6, V0eiu6, C1eiu6, J1eiu6, Q1eiu6, X1eiu6, E2eiu6, L2eiu6;
wire S2eiu6, Z2eiu6, G3eiu6, N3eiu6, U3eiu6, B4eiu6, I4eiu6, P4eiu6, W4eiu6, D5eiu6;
wire K5eiu6, R5eiu6, Y5eiu6, F6eiu6, M6eiu6, T6eiu6, A7eiu6, H7eiu6, O7eiu6, V7eiu6;
wire C8eiu6, J8eiu6, Q8eiu6, X8eiu6, E9eiu6, L9eiu6, S9eiu6, Z9eiu6, Gaeiu6, Naeiu6;
wire Uaeiu6, Bbeiu6, Ibeiu6, Pbeiu6, Wbeiu6, Dceiu6, Kceiu6, Rceiu6, Yceiu6, Fdeiu6;
wire Mdeiu6, Tdeiu6, Aeeiu6, Heeiu6, Oeeiu6, Veeiu6, Cfeiu6, Jfeiu6, Qfeiu6, Xfeiu6;
wire Egeiu6, Lgeiu6, Sgeiu6, Zgeiu6, Gheiu6, Nheiu6, Uheiu6, Bieiu6, Iieiu6, Pieiu6;
wire Wieiu6, Djeiu6, Kjeiu6, Rjeiu6, Yjeiu6, Fkeiu6, Mkeiu6, Tkeiu6, Aleiu6, Hleiu6;
wire Oleiu6, Vleiu6, Cmeiu6, Jmeiu6, Qmeiu6, Xmeiu6, Eneiu6, Lneiu6, Sneiu6, Zneiu6;
wire Goeiu6, Noeiu6, Uoeiu6, Bpeiu6, Ipeiu6, Ppeiu6, Wpeiu6, Dqeiu6, Kqeiu6, Rqeiu6;
wire Yqeiu6, Freiu6, Mreiu6, Treiu6, Aseiu6, Hseiu6, Oseiu6, Vseiu6, Cteiu6, Jteiu6;
wire Qteiu6, Xteiu6, Eueiu6, Lueiu6, Sueiu6, Zueiu6, Gveiu6, Nveiu6, Uveiu6, Bweiu6;
wire Iweiu6, Pweiu6, Wweiu6, Dxeiu6, Kxeiu6, Rxeiu6, Yxeiu6, Fyeiu6, Myeiu6, Tyeiu6;
wire Azeiu6, Hzeiu6, Ozeiu6, Vzeiu6, C0fiu6, J0fiu6, Q0fiu6, X0fiu6, E1fiu6, L1fiu6;
wire S1fiu6, Z1fiu6, G2fiu6, N2fiu6, U2fiu6, B3fiu6, I3fiu6, P3fiu6, W3fiu6, D4fiu6;
wire K4fiu6, R4fiu6, Y4fiu6, F5fiu6, M5fiu6, T5fiu6, A6fiu6, H6fiu6, O6fiu6, V6fiu6;
wire C7fiu6, J7fiu6, Q7fiu6, X7fiu6, E8fiu6, L8fiu6, S8fiu6, Z8fiu6, G9fiu6, N9fiu6;
wire U9fiu6, Bafiu6, Iafiu6, Pafiu6, Wafiu6, Dbfiu6, Kbfiu6, Rbfiu6, Ybfiu6, Fcfiu6;
wire Mcfiu6, Tcfiu6, Adfiu6, Hdfiu6, Odfiu6, Vdfiu6, Cefiu6, Jefiu6, Qefiu6, Xefiu6;
wire Effiu6, Lffiu6, Sffiu6, Zffiu6, Ggfiu6, Ngfiu6, Ugfiu6, Bhfiu6, Ihfiu6, Phfiu6;
wire Whfiu6, Difiu6, Kifiu6, Rifiu6, Yifiu6, Fjfiu6, Mjfiu6, Tjfiu6, Akfiu6, Hkfiu6;
wire Okfiu6, Vkfiu6, Clfiu6, Jlfiu6, Qlfiu6, Xlfiu6, Emfiu6, Lmfiu6, Smfiu6, Zmfiu6;
wire Gnfiu6, Nnfiu6, Unfiu6, Bofiu6, Iofiu6, Pofiu6, Wofiu6, Dpfiu6, Kpfiu6, Rpfiu6;
wire Ypfiu6, Fqfiu6, Mqfiu6, Tqfiu6, Arfiu6, Hrfiu6, Orfiu6, Vrfiu6, Csfiu6, Jsfiu6;
wire Qsfiu6, Xsfiu6, Etfiu6, Ltfiu6, Stfiu6, Ztfiu6, Gufiu6, Nufiu6, Uufiu6, Bvfiu6;
wire Ivfiu6, Pvfiu6, Wvfiu6, Dwfiu6, Kwfiu6, Rwfiu6, Ywfiu6, Fxfiu6, Mxfiu6, Txfiu6;
wire Ayfiu6, Hyfiu6, Oyfiu6, Vyfiu6, Czfiu6, Jzfiu6, Qzfiu6, Xzfiu6, E0giu6, L0giu6;
wire S0giu6, Z0giu6, G1giu6, N1giu6, U1giu6, B2giu6, I2giu6, P2giu6, W2giu6, D3giu6;
wire K3giu6, R3giu6, Y3giu6, F4giu6, M4giu6, T4giu6, A5giu6, H5giu6, O5giu6, V5giu6;
wire C6giu6, J6giu6, Q6giu6, X6giu6, E7giu6, L7giu6, S7giu6, Z7giu6, G8giu6, N8giu6;
wire U8giu6, B9giu6, I9giu6, P9giu6, W9giu6, Dagiu6, Kagiu6, Ragiu6, Yagiu6, Fbgiu6;
wire Mbgiu6, Tbgiu6, Acgiu6, Hcgiu6, Ocgiu6, Vcgiu6, Cdgiu6, Jdgiu6, Qdgiu6, Xdgiu6;
wire Eegiu6, Legiu6, Segiu6, Zegiu6, Gfgiu6, Nfgiu6, Ufgiu6, Bggiu6, Iggiu6, Pggiu6;
wire Wggiu6, Dhgiu6, Khgiu6, Rhgiu6, Yhgiu6, Figiu6, Migiu6, Tigiu6, Ajgiu6, Hjgiu6;
wire Ojgiu6, Vjgiu6, Ckgiu6, Jkgiu6, Qkgiu6, Xkgiu6, Elgiu6, Llgiu6, Slgiu6, Zlgiu6;
wire Gmgiu6, Nmgiu6, Umgiu6, Bngiu6, Ingiu6, Pngiu6, Wngiu6, Dogiu6, Kogiu6, Rogiu6;
wire Yogiu6, Fpgiu6, Mpgiu6, Tpgiu6, Aqgiu6, Hqgiu6, Oqgiu6, Vqgiu6, Crgiu6, Jrgiu6;
wire Qrgiu6, Xrgiu6, Esgiu6, Lsgiu6, Ssgiu6, Zsgiu6, Gtgiu6, Ntgiu6, Utgiu6, Bugiu6;
wire Iugiu6, Pugiu6, Wugiu6, Dvgiu6, Kvgiu6, Rvgiu6, Yvgiu6, Fwgiu6, Mwgiu6, Twgiu6;
wire Axgiu6, Hxgiu6, Oxgiu6, Vxgiu6, Cygiu6, Jygiu6, Qygiu6, Xygiu6, Ezgiu6, Lzgiu6;
wire Szgiu6, Zzgiu6, G0hiu6, N0hiu6, U0hiu6, B1hiu6, I1hiu6, P1hiu6, W1hiu6, D2hiu6;
wire K2hiu6, R2hiu6, Y2hiu6, F3hiu6, M3hiu6, T3hiu6, A4hiu6, H4hiu6, O4hiu6, V4hiu6;
wire C5hiu6, J5hiu6, Q5hiu6, X5hiu6, E6hiu6, L6hiu6, S6hiu6, Z6hiu6, G7hiu6, N7hiu6;
wire U7hiu6, B8hiu6, I8hiu6, P8hiu6, W8hiu6, D9hiu6, K9hiu6, R9hiu6, Y9hiu6, Fahiu6;
wire Mahiu6, Tahiu6, Abhiu6, Hbhiu6, Obhiu6, Vbhiu6, Cchiu6, Jchiu6, Qchiu6, Xchiu6;
wire Edhiu6, Ldhiu6, Sdhiu6, Zdhiu6, Gehiu6, Nehiu6, Uehiu6, Bfhiu6, Ifhiu6, Pfhiu6;
wire Wfhiu6, Dghiu6, Kghiu6, Rghiu6, Yghiu6, Fhhiu6, Mhhiu6, Thhiu6, Aihiu6, Hihiu6;
wire Oihiu6, Vihiu6, Cjhiu6, Jjhiu6, Qjhiu6, Xjhiu6, Ekhiu6, Lkhiu6, Skhiu6, Zkhiu6;
wire Glhiu6, Nlhiu6, Ulhiu6, Bmhiu6, Imhiu6, Pmhiu6, Wmhiu6, Dnhiu6, Knhiu6, Rnhiu6;
wire Ynhiu6, Fohiu6, Mohiu6, Tohiu6, Aphiu6, Hphiu6, Ophiu6, Vphiu6, Cqhiu6, Jqhiu6;
wire Qqhiu6, Xqhiu6, Erhiu6, Lrhiu6, Srhiu6, Zrhiu6, Gshiu6, Nshiu6, Ushiu6, Bthiu6;
wire Ithiu6, Pthiu6, Wthiu6, Duhiu6, Kuhiu6, Ruhiu6, Yuhiu6, Fvhiu6, Mvhiu6, Tvhiu6;
wire Awhiu6, Hwhiu6, Owhiu6, Vwhiu6, Cxhiu6, Jxhiu6, Qxhiu6, Xxhiu6, Eyhiu6, Lyhiu6;
wire Syhiu6, Zyhiu6, Gzhiu6, Nzhiu6, Uzhiu6, B0iiu6, I0iiu6, P0iiu6, W0iiu6, D1iiu6;
wire K1iiu6, R1iiu6, Y1iiu6, F2iiu6, M2iiu6, T2iiu6, A3iiu6, H3iiu6, O3iiu6, V3iiu6;
wire C4iiu6, J4iiu6, Q4iiu6, X4iiu6, E5iiu6, L5iiu6, S5iiu6, Z5iiu6, G6iiu6, N6iiu6;
wire U6iiu6, B7iiu6, I7iiu6, P7iiu6, W7iiu6, D8iiu6, K8iiu6, R8iiu6, Y8iiu6, F9iiu6;
wire M9iiu6, T9iiu6, Aaiiu6, Haiiu6, Oaiiu6, Vaiiu6, Cbiiu6, Jbiiu6, Qbiiu6, Xbiiu6;
wire Eciiu6, Lciiu6, Sciiu6, Zciiu6, Gdiiu6, Ndiiu6, Udiiu6, Beiiu6, Ieiiu6, Peiiu6;
wire Weiiu6, Dfiiu6, Kfiiu6, Rfiiu6, Yfiiu6, Fgiiu6, Mgiiu6, Tgiiu6, Ahiiu6, Hhiiu6;
wire Ohiiu6, Vhiiu6, Ciiiu6, Jiiiu6, Qiiiu6, Xiiiu6, Ejiiu6, Ljiiu6, Sjiiu6, Zjiiu6;
wire Gkiiu6, Nkiiu6, Ukiiu6, Bliiu6, Iliiu6, Pliiu6, Wliiu6, Dmiiu6, Kmiiu6, Rmiiu6;
wire Ymiiu6, Fniiu6, Mniiu6, Tniiu6, Aoiiu6, Hoiiu6, Ooiiu6, Voiiu6, Cpiiu6, Jpiiu6;
wire Qpiiu6, Xpiiu6, Eqiiu6, Lqiiu6, Sqiiu6, Zqiiu6, Griiu6, Nriiu6, Uriiu6, Bsiiu6;
wire Isiiu6, Psiiu6, Wsiiu6, Dtiiu6, Ktiiu6, Rtiiu6, Ytiiu6, Fuiiu6, Muiiu6, Tuiiu6;
wire Aviiu6, Hviiu6, Oviiu6, Vviiu6, Cwiiu6, Jwiiu6, Qwiiu6, Xwiiu6, Exiiu6, Lxiiu6;
wire Sxiiu6, Zxiiu6, Gyiiu6, Nyiiu6, Uyiiu6, Bziiu6, Iziiu6, Pziiu6, Wziiu6, D0jiu6;
wire K0jiu6, R0jiu6, Y0jiu6, F1jiu6, M1jiu6, T1jiu6, A2jiu6, H2jiu6, O2jiu6, V2jiu6;
wire C3jiu6, J3jiu6, Q3jiu6, X3jiu6, E4jiu6, L4jiu6, S4jiu6, Z4jiu6, G5jiu6, N5jiu6;
wire U5jiu6, B6jiu6, I6jiu6, P6jiu6, W6jiu6, D7jiu6, K7jiu6, R7jiu6, Y7jiu6, F8jiu6;
wire M8jiu6, T8jiu6, A9jiu6, H9jiu6, O9jiu6, V9jiu6, Cajiu6, Jajiu6, Qajiu6, Xajiu6;
wire Ebjiu6, Lbjiu6, Sbjiu6, Zbjiu6, Gcjiu6, Ncjiu6, Ucjiu6, Bdjiu6, Idjiu6, Pdjiu6;
wire Wdjiu6, Dejiu6, Kejiu6, Rejiu6, Yejiu6, Ffjiu6, Mfjiu6, Tfjiu6, Agjiu6, Hgjiu6;
wire Ogjiu6, Vgjiu6, Chjiu6, Jhjiu6, Qhjiu6, Xhjiu6, Eijiu6, Lijiu6, Sijiu6, Zijiu6;
wire Gjjiu6, Njjiu6, Ujjiu6, Bkjiu6, Ikjiu6, Pkjiu6, Wkjiu6, Dljiu6, Kljiu6, Rljiu6;
wire Yljiu6, Fmjiu6, Mmjiu6, Tmjiu6, Anjiu6, Hnjiu6, Onjiu6, Vnjiu6, Cojiu6, Jojiu6;
wire Qojiu6, Xojiu6, Epjiu6, Lpjiu6, Spjiu6, Zpjiu6, Gqjiu6, Nqjiu6, Uqjiu6, Brjiu6;
wire Irjiu6, Prjiu6, Wrjiu6, Dsjiu6, Ksjiu6, Rsjiu6, Ysjiu6, Ftjiu6, Mtjiu6, Ttjiu6;
wire Aujiu6, Hujiu6, Oujiu6, Vujiu6, Cvjiu6, Jvjiu6, Qvjiu6, Xvjiu6, Ewjiu6, Lwjiu6;
wire Swjiu6, Zwjiu6, Gxjiu6, Nxjiu6, Uxjiu6, Byjiu6, Iyjiu6, Pyjiu6, Wyjiu6, Dzjiu6;
wire Kzjiu6, Rzjiu6, Yzjiu6, F0kiu6, M0kiu6, T0kiu6, A1kiu6, H1kiu6, O1kiu6, V1kiu6;
wire C2kiu6, J2kiu6, Q2kiu6, X2kiu6, E3kiu6, L3kiu6, S3kiu6, Z3kiu6, G4kiu6, N4kiu6;
wire U4kiu6, B5kiu6, I5kiu6, P5kiu6, W5kiu6, D6kiu6, K6kiu6, R6kiu6, Y6kiu6, F7kiu6;
wire M7kiu6, T7kiu6, A8kiu6, H8kiu6, O8kiu6, V8kiu6, C9kiu6, J9kiu6, Q9kiu6, X9kiu6;
wire Eakiu6, Lakiu6, Sakiu6, Zakiu6, Gbkiu6, Nbkiu6, Ubkiu6, Bckiu6, Ickiu6, Pckiu6;
wire Wckiu6, Ddkiu6, Kdkiu6, Rdkiu6, Ydkiu6, Fekiu6, Mekiu6, Tekiu6, Afkiu6, Hfkiu6;
wire Ofkiu6, Vfkiu6, Cgkiu6, Jgkiu6, Qgkiu6, Xgkiu6, Ehkiu6, Lhkiu6, Shkiu6, Zhkiu6;
wire Gikiu6, Nikiu6, Uikiu6, Bjkiu6, Ijkiu6, Pjkiu6, Wjkiu6, Dkkiu6, Kkkiu6, Rkkiu6;
wire Ykkiu6, Flkiu6, Mlkiu6, Tlkiu6, Amkiu6, Hmkiu6, Omkiu6, Vmkiu6, Cnkiu6, Jnkiu6;
wire Qnkiu6, Xnkiu6, Eokiu6, Lokiu6, Sokiu6, Zokiu6, Gpkiu6, Npkiu6, Upkiu6, Bqkiu6;
wire Iqkiu6, Pqkiu6, Wqkiu6, Drkiu6, Krkiu6, Rrkiu6, Yrkiu6, Fskiu6, Mskiu6, Tskiu6;
wire Atkiu6, Htkiu6, Otkiu6, Vtkiu6, Cukiu6, Jukiu6, Qukiu6, Xukiu6, Evkiu6, Lvkiu6;
wire Svkiu6, Zvkiu6, Gwkiu6, Nwkiu6, Uwkiu6, Bxkiu6, Ixkiu6, Pxkiu6, Wxkiu6, Dykiu6;
wire Kykiu6, Rykiu6, Yykiu6, Fzkiu6, Mzkiu6, Tzkiu6, A0liu6, H0liu6, O0liu6, V0liu6;
wire C1liu6, J1liu6, Q1liu6, X1liu6, E2liu6, L2liu6, S2liu6, Z2liu6, G3liu6, N3liu6;
wire U3liu6, B4liu6, I4liu6, P4liu6, W4liu6, D5liu6, K5liu6, R5liu6, Y5liu6, F6liu6;
wire M6liu6, T6liu6, A7liu6, H7liu6, O7liu6, V7liu6, C8liu6, J8liu6, Q8liu6, X8liu6;
wire E9liu6, L9liu6, S9liu6, Z9liu6, Galiu6, Naliu6, Ualiu6, Bbliu6, Ibliu6, Pbliu6;
wire Wbliu6, Dcliu6, Kcliu6, Rcliu6, Ycliu6, Fdliu6, Mdliu6, Tdliu6, Aeliu6, Heliu6;
wire Oeliu6, Veliu6, Cfliu6, Jfliu6, Qfliu6, Xfliu6, Egliu6, Lgliu6, Sgliu6, Zgliu6;
wire Ghliu6, Nhliu6, Uhliu6, Biliu6, Iiliu6, Piliu6, Wiliu6, Djliu6, Kjliu6, Rjliu6;
wire Yjliu6, Fkliu6, Mkliu6, Tkliu6, Alliu6, Hlliu6, Olliu6, Vlliu6, Cmliu6, Jmliu6;
wire Qmliu6, Xmliu6, Enliu6, Lnliu6, Snliu6, Znliu6, Goliu6, Noliu6, Uoliu6, Bpliu6;
wire Ipliu6, Ppliu6, Wpliu6, Dqliu6, Kqliu6, Rqliu6, Yqliu6, Frliu6, Mrliu6, Trliu6;
wire Asliu6, Hsliu6, Osliu6, Vsliu6, Ctliu6, Jtliu6, Qtliu6, Xtliu6, Euliu6, Luliu6;
wire Suliu6, Zuliu6, Gvliu6, Nvliu6, Uvliu6, Bwliu6, Iwliu6, Pwliu6, Wwliu6, Dxliu6;
wire Kxliu6, Rxliu6, Yxliu6, Fyliu6, Myliu6, Tyliu6, Azliu6, Hzliu6, Ozliu6, Vzliu6;
wire C0miu6, J0miu6, Q0miu6, X0miu6, E1miu6, L1miu6, S1miu6, Z1miu6, G2miu6, N2miu6;
wire U2miu6, B3miu6, I3miu6, P3miu6, W3miu6, D4miu6, K4miu6, R4miu6, Y4miu6, F5miu6;
wire M5miu6, T5miu6, A6miu6, H6miu6, O6miu6, V6miu6, C7miu6, J7miu6, Q7miu6, X7miu6;
wire E8miu6, L8miu6, S8miu6, Z8miu6, G9miu6, N9miu6, U9miu6, Bamiu6, Iamiu6, Pamiu6;
wire Wamiu6, Dbmiu6, Kbmiu6, Rbmiu6, Ybmiu6, Fcmiu6, Mcmiu6, Tcmiu6, Admiu6, Hdmiu6;
wire Odmiu6, Vdmiu6, Cemiu6, Jemiu6, Qemiu6, Xemiu6, Efmiu6, Lfmiu6, Sfmiu6, Zfmiu6;
wire Ggmiu6, Ngmiu6, Ugmiu6, Bhmiu6, Ihmiu6, Phmiu6, Whmiu6, Dimiu6, Kimiu6, Rimiu6;
wire Yimiu6, Fjmiu6, Mjmiu6, Tjmiu6, Akmiu6, Hkmiu6, Okmiu6, Vkmiu6, Clmiu6, Jlmiu6;
wire Qlmiu6, Xlmiu6, Emmiu6, Lmmiu6, Smmiu6, Zmmiu6, Gnmiu6, Nnmiu6, Unmiu6, Bomiu6;
wire Iomiu6, Pomiu6, Womiu6, Dpmiu6, Kpmiu6, Rpmiu6, Ypmiu6, Fqmiu6, Mqmiu6, Tqmiu6;
wire Armiu6, Hrmiu6, Ormiu6, Vrmiu6, Csmiu6, Jsmiu6, Qsmiu6, Xsmiu6, Etmiu6, Ltmiu6;
wire Stmiu6, Ztmiu6, Gumiu6, Numiu6, Uumiu6, Bvmiu6, Ivmiu6, Pvmiu6, Wvmiu6, Dwmiu6;
wire Kwmiu6, Rwmiu6, Ywmiu6, Fxmiu6, Mxmiu6, Txmiu6, Aymiu6, Hymiu6, Oymiu6, Vymiu6;
wire Czmiu6, Jzmiu6, Qzmiu6, Xzmiu6, E0niu6, L0niu6, S0niu6, Z0niu6, G1niu6, N1niu6;
wire U1niu6, B2niu6, I2niu6, P2niu6, W2niu6, D3niu6, K3niu6, R3niu6, Y3niu6, F4niu6;
wire M4niu6, T4niu6, A5niu6, H5niu6, O5niu6, V5niu6, C6niu6, J6niu6, Q6niu6, X6niu6;
wire E7niu6, L7niu6, S7niu6, Z7niu6, G8niu6, N8niu6, U8niu6, B9niu6, I9niu6, P9niu6;
wire W9niu6, Daniu6, Kaniu6, Raniu6, Yaniu6, Fbniu6, Mbniu6, Tbniu6, Acniu6, Hcniu6;
wire Ocniu6, Vcniu6, Cdniu6, Jdniu6, Qdniu6, Xdniu6, Eeniu6, Leniu6, Seniu6, Zeniu6;
wire Gfniu6, Nfniu6, Ufniu6, Bgniu6, Igniu6, Pgniu6, Wgniu6, Dhniu6, Khniu6, Rhniu6;
wire Yhniu6, Finiu6, Miniu6, Tiniu6, Ajniu6, Hjniu6, Ojniu6, Vjniu6, Ckniu6, Jkniu6;
wire Qkniu6, Xkniu6, Elniu6, Llniu6, Slniu6, Zlniu6, Gmniu6, Nmniu6, Umniu6, Bnniu6;
wire Inniu6, Pnniu6, Wnniu6, Doniu6, Koniu6, Roniu6, Yoniu6, Fpniu6, Mpniu6, Tpniu6;
wire Aqniu6, Hqniu6, Oqniu6, Vqniu6, Crniu6, Jrniu6, Qrniu6, Xrniu6, Esniu6, Lsniu6;
wire Ssniu6, Zsniu6, Gtniu6, Ntniu6, Utniu6, Buniu6, Iuniu6, Puniu6, Wuniu6, Dvniu6;
wire Kvniu6, Rvniu6, Yvniu6, Fwniu6, Mwniu6, Twniu6, Axniu6, Hxniu6, Oxniu6, Vxniu6;
wire Cyniu6, Jyniu6, Qyniu6, Xyniu6, Ezniu6, Lzniu6, Szniu6, Zzniu6, G0oiu6, N0oiu6;
wire U0oiu6, B1oiu6, I1oiu6, P1oiu6, W1oiu6, D2oiu6, K2oiu6, R2oiu6, Y2oiu6, F3oiu6;
wire M3oiu6, T3oiu6, A4oiu6, H4oiu6, O4oiu6, V4oiu6, C5oiu6, J5oiu6, Q5oiu6, X5oiu6;
wire E6oiu6, L6oiu6, S6oiu6, Z6oiu6, G7oiu6, N7oiu6, U7oiu6, B8oiu6, I8oiu6, P8oiu6;
wire W8oiu6, D9oiu6, K9oiu6, R9oiu6, Y9oiu6, Faoiu6, Maoiu6, Taoiu6, Aboiu6, Hboiu6;
wire Oboiu6, Vboiu6, Ccoiu6, Jcoiu6, Qcoiu6, Xcoiu6, Edoiu6, Ldoiu6, Sdoiu6, Zdoiu6;
wire Geoiu6, Neoiu6, Ueoiu6, Bfoiu6, Ifoiu6, Pfoiu6, Wfoiu6, Dgoiu6, Kgoiu6, Rgoiu6;
wire Ygoiu6, Fhoiu6, Mhoiu6, Thoiu6, Aioiu6, Hioiu6, Oioiu6, Vioiu6, Cjoiu6, Jjoiu6;
wire Qjoiu6, Xjoiu6, Ekoiu6, Lkoiu6, Skoiu6, Zkoiu6, Gloiu6, Nloiu6, Uloiu6, Bmoiu6;
wire Imoiu6, Pmoiu6, Wmoiu6, Dnoiu6, Knoiu6, Rnoiu6, Ynoiu6, Fooiu6, Mooiu6, Tooiu6;
wire Apoiu6, Hpoiu6, Opoiu6, Vpoiu6, Cqoiu6, Jqoiu6, Qqoiu6, Xqoiu6, Eroiu6, Lroiu6;
wire Sroiu6, Zroiu6, Gsoiu6, Nsoiu6, Usoiu6, Btoiu6, Itoiu6, Ptoiu6, Wtoiu6, Duoiu6;
wire Kuoiu6, Ruoiu6, Yuoiu6, Fvoiu6, Mvoiu6, Tvoiu6, Awoiu6, Hwoiu6, Owoiu6, Vwoiu6;
wire Cxoiu6, Jxoiu6, Qxoiu6, Xxoiu6, Eyoiu6, Lyoiu6, Syoiu6, Zyoiu6, Gzoiu6, Nzoiu6;
wire Uzoiu6, B0piu6, I0piu6, P0piu6, W0piu6, D1piu6, K1piu6, R1piu6, Y1piu6, F2piu6;
wire M2piu6, T2piu6, A3piu6, H3piu6, O3piu6, V3piu6, C4piu6, J4piu6, Q4piu6, X4piu6;
wire E5piu6, L5piu6, S5piu6, Z5piu6, G6piu6, N6piu6, U6piu6, B7piu6, I7piu6, P7piu6;
wire W7piu6, D8piu6, K8piu6, R8piu6, Y8piu6, F9piu6, M9piu6, T9piu6, Aapiu6, Hapiu6;
wire Oapiu6, Vapiu6, Cbpiu6, Jbpiu6, Qbpiu6, Xbpiu6, Ecpiu6, Lcpiu6, Scpiu6, Zcpiu6;
wire Gdpiu6, Ndpiu6, Udpiu6, Bepiu6, Iepiu6, Pepiu6, Wepiu6, Dfpiu6, Kfpiu6, Rfpiu6;
wire Yfpiu6, Fgpiu6, Mgpiu6, Tgpiu6, Ahpiu6, Hhpiu6, Ohpiu6, Vhpiu6, Cipiu6, Jipiu6;
wire Qipiu6, Xipiu6, Ejpiu6, Ljpiu6, Sjpiu6, Zjpiu6, Gkpiu6, Nkpiu6, Ukpiu6, Blpiu6;
wire Ilpiu6, Plpiu6, Wlpiu6, Dmpiu6, Kmpiu6, Rmpiu6, Ympiu6, Fnpiu6, Mnpiu6, Tnpiu6;
wire Aopiu6, Hopiu6, Oopiu6, Vopiu6, Cppiu6, Jppiu6, Qppiu6, Xppiu6, Eqpiu6, Lqpiu6;
wire Sqpiu6, Zqpiu6, Grpiu6, Nrpiu6, Urpiu6, Bspiu6, Ispiu6, Pspiu6, Wspiu6, Dtpiu6;
wire Ktpiu6, Rtpiu6, Ytpiu6, Fupiu6, Mupiu6, Tupiu6, Avpiu6, Hvpiu6, Ovpiu6, Vvpiu6;
wire Cwpiu6, Jwpiu6, Qwpiu6, Xwpiu6, Expiu6, Lxpiu6, Sxpiu6, Zxpiu6, Gypiu6, Nypiu6;
wire Uypiu6, Bzpiu6, Izpiu6, Pzpiu6, Wzpiu6, D0qiu6, K0qiu6, R0qiu6, Y0qiu6, F1qiu6;
wire M1qiu6, T1qiu6, A2qiu6, H2qiu6, O2qiu6, V2qiu6, C3qiu6, J3qiu6, Q3qiu6, X3qiu6;
wire E4qiu6, L4qiu6, S4qiu6, Z4qiu6, G5qiu6, N5qiu6, U5qiu6, B6qiu6, I6qiu6, P6qiu6;
wire W6qiu6, D7qiu6, K7qiu6, R7qiu6, Y7qiu6, F8qiu6, M8qiu6, T8qiu6, A9qiu6, H9qiu6;
wire O9qiu6, V9qiu6, Caqiu6, Jaqiu6, Qaqiu6, Xaqiu6, Ebqiu6, Lbqiu6, Sbqiu6, Zbqiu6;
wire Gcqiu6, Ncqiu6, Ucqiu6, Bdqiu6, Idqiu6, Pdqiu6, Wdqiu6, Deqiu6, Keqiu6, Reqiu6;
wire Yeqiu6, Ffqiu6, Mfqiu6, Tfqiu6, Agqiu6, Hgqiu6, Ogqiu6, Vgqiu6, Chqiu6, Jhqiu6;
wire Qhqiu6, Xhqiu6, Eiqiu6, Liqiu6, Siqiu6, Ziqiu6, Gjqiu6, Njqiu6, Ujqiu6, Bkqiu6;
wire Ikqiu6, Pkqiu6, Wkqiu6, Dlqiu6, Klqiu6, Rlqiu6, Ylqiu6, Fmqiu6, Mmqiu6, Tmqiu6;
wire Anqiu6, Hnqiu6, Onqiu6, Vnqiu6, Coqiu6, Joqiu6, Qoqiu6, Xoqiu6, Epqiu6, Lpqiu6;
wire Spqiu6, Zpqiu6, Gqqiu6, Nqqiu6, Uqqiu6, Brqiu6, Irqiu6, Prqiu6, Wrqiu6, Dsqiu6;
wire Ksqiu6, Rsqiu6, Ysqiu6, Ftqiu6, Mtqiu6, Ttqiu6, Auqiu6, Huqiu6, Ouqiu6, Vuqiu6;
wire Cvqiu6, Jvqiu6, Qvqiu6, Xvqiu6, Ewqiu6, Lwqiu6, Swqiu6, Zwqiu6, Gxqiu6, Nxqiu6;
wire Uxqiu6, Byqiu6, Iyqiu6, Pyqiu6, Wyqiu6, Dzqiu6, Kzqiu6, Rzqiu6, Yzqiu6, F0riu6;
wire M0riu6, T0riu6, A1riu6, H1riu6, O1riu6, V1riu6, C2riu6, J2riu6, Q2riu6, X2riu6;
wire E3riu6, L3riu6, S3riu6, Z3riu6, G4riu6, N4riu6, U4riu6, B5riu6, I5riu6, P5riu6;
wire W5riu6, D6riu6, K6riu6, R6riu6, Y6riu6, F7riu6, M7riu6, T7riu6, A8riu6, H8riu6;
wire O8riu6, V8riu6, C9riu6, J9riu6, Q9riu6, X9riu6, Eariu6, Lariu6, Sariu6, Zariu6;
wire Gbriu6, Nbriu6, Ubriu6, Bcriu6, Icriu6, Pcriu6, Wcriu6, Ddriu6, Kdriu6, Rdriu6;
wire Ydriu6, Feriu6, Meriu6, Teriu6, Afriu6, Hfriu6, Ofriu6, Vfriu6, Cgriu6, Jgriu6;
wire Qgriu6, Xgriu6, Ehriu6, Lhriu6, Shriu6, Zhriu6, Giriu6, Niriu6, Uiriu6, Bjriu6;
wire Ijriu6, Pjriu6, Wjriu6, Dkriu6, Kkriu6, Rkriu6, Ykriu6, Flriu6, Mlriu6, Tlriu6;
wire Amriu6, Hmriu6, Omriu6, Vmriu6, Cnriu6, Jnriu6, Qnriu6, Xnriu6, Eoriu6, Loriu6;
wire Soriu6, Zoriu6, Gpriu6, Npriu6, Upriu6, Bqriu6, Iqriu6, Pqriu6, Wqriu6, Drriu6;
wire Krriu6, Rrriu6, Yrriu6, Fsriu6, Msriu6, Tsriu6, Atriu6, Htriu6, Otriu6, Vtriu6;
wire Curiu6, Juriu6, Quriu6, Xuriu6, Evriu6, Lvriu6, Svriu6, Zvriu6, Gwriu6, Nwriu6;
wire Uwriu6, Bxriu6, Ixriu6, Pxriu6, Wxriu6, Dyriu6, Kyriu6, Ryriu6, Yyriu6, Fzriu6;
wire Mzriu6, Tzriu6, A0siu6, H0siu6, O0siu6, V0siu6, C1siu6, J1siu6, Q1siu6, X1siu6;
wire E2siu6, L2siu6, S2siu6, Z2siu6, G3siu6, N3siu6, U3siu6, B4siu6, I4siu6, P4siu6;
wire W4siu6, D5siu6, K5siu6, R5siu6, Y5siu6, F6siu6, M6siu6, T6siu6, A7siu6, H7siu6;
wire O7siu6, V7siu6, C8siu6, J8siu6, Q8siu6, X8siu6, E9siu6, L9siu6, S9siu6, Z9siu6;
wire Gasiu6, Nasiu6, Uasiu6, Bbsiu6, Ibsiu6, Pbsiu6, Wbsiu6, Dcsiu6, Kcsiu6, Rcsiu6;
wire Ycsiu6, Fdsiu6, Mdsiu6, Tdsiu6, Aesiu6, Hesiu6, Oesiu6, Vesiu6, Cfsiu6, Jfsiu6;
wire Qfsiu6, Xfsiu6, Egsiu6, Lgsiu6, Sgsiu6, Zgsiu6, Ghsiu6, Nhsiu6, Uhsiu6, Bisiu6;
wire Iisiu6, Pisiu6, Wisiu6, Djsiu6, Kjsiu6, Rjsiu6, Yjsiu6, Fksiu6, Mksiu6, Tksiu6;
wire Alsiu6, Hlsiu6, Olsiu6, Vlsiu6, Cmsiu6, Jmsiu6, Qmsiu6, Xmsiu6, Ensiu6, Lnsiu6;
wire Snsiu6, Znsiu6, Gosiu6, Nosiu6, Uosiu6, Bpsiu6, Ipsiu6, Ppsiu6, Wpsiu6, Dqsiu6;
wire Kqsiu6, Rqsiu6, Yqsiu6, Frsiu6, Mrsiu6, Trsiu6, Assiu6, Hssiu6, Ossiu6, Vssiu6;
wire Ctsiu6, Jtsiu6, Qtsiu6, Xtsiu6, Eusiu6, Lusiu6, Susiu6, Zusiu6, Gvsiu6, Nvsiu6;
wire Uvsiu6, Bwsiu6, Iwsiu6, Pwsiu6, Wwsiu6, Dxsiu6, Kxsiu6, Rxsiu6, Yxsiu6, Fysiu6;
wire Mysiu6, Tysiu6, Azsiu6, Hzsiu6, Ozsiu6, Vzsiu6, C0tiu6, J0tiu6, Q0tiu6, X0tiu6;
wire E1tiu6, L1tiu6, S1tiu6, Z1tiu6, G2tiu6, N2tiu6, U2tiu6, B3tiu6, I3tiu6, P3tiu6;
wire W3tiu6, D4tiu6, K4tiu6, R4tiu6, Y4tiu6, F5tiu6, M5tiu6, T5tiu6, A6tiu6, H6tiu6;
wire O6tiu6, V6tiu6, C7tiu6, J7tiu6, Q7tiu6, X7tiu6, E8tiu6, L8tiu6, S8tiu6, Z8tiu6;
wire G9tiu6, N9tiu6, U9tiu6, Batiu6, Iatiu6, Patiu6, Watiu6, Dbtiu6, Kbtiu6, Rbtiu6;
wire Ybtiu6, Fctiu6, Mctiu6, Tctiu6, Adtiu6, Hdtiu6, Odtiu6, Vdtiu6, Cetiu6, Jetiu6;
wire Qetiu6, Xetiu6, Eftiu6, Lftiu6, Sftiu6, Zftiu6, Ggtiu6, Ngtiu6, Ugtiu6, Bhtiu6;
wire Ihtiu6, Phtiu6, Whtiu6, Ditiu6, Kitiu6, Ritiu6, Yitiu6, Fjtiu6, Mjtiu6, Tjtiu6;
wire Aktiu6, Hktiu6, Oktiu6, Vktiu6, Cltiu6, Jltiu6, Qltiu6, Xltiu6, Emtiu6, Lmtiu6;
wire Smtiu6, Zmtiu6, Gntiu6, Nntiu6, Untiu6, Botiu6, Iotiu6, Potiu6, Wotiu6, Dptiu6;
wire Kptiu6, Rptiu6, Yptiu6, Fqtiu6, Mqtiu6, Tqtiu6, Artiu6, Hrtiu6, Ortiu6, Vrtiu6;
wire Cstiu6, Jstiu6, Qstiu6, Xstiu6, Ettiu6, Lttiu6, Sttiu6, Zttiu6, Gutiu6, Nutiu6;
wire Uutiu6, Bvtiu6, Ivtiu6, Pvtiu6, Wvtiu6, Dwtiu6, Kwtiu6, Rwtiu6, Ywtiu6, Fxtiu6;
wire Mxtiu6, Txtiu6, Aytiu6, Hytiu6, Oytiu6, Vytiu6, Cztiu6, Jztiu6, Qztiu6, Xztiu6;
wire E0uiu6, L0uiu6, S0uiu6, Z0uiu6, G1uiu6, N1uiu6, U1uiu6, B2uiu6, I2uiu6, P2uiu6;
wire W2uiu6, D3uiu6, K3uiu6, R3uiu6, Y3uiu6, F4uiu6, M4uiu6, T4uiu6, A5uiu6, H5uiu6;
wire O5uiu6, V5uiu6, C6uiu6, J6uiu6, Q6uiu6, X6uiu6, E7uiu6, L7uiu6, S7uiu6, Z7uiu6;
wire G8uiu6, N8uiu6, U8uiu6, B9uiu6, I9uiu6, P9uiu6, W9uiu6, Dauiu6, Kauiu6, Rauiu6;
wire Yauiu6, Fbuiu6, Mbuiu6, Tbuiu6, Acuiu6, Hcuiu6, Ocuiu6, Vcuiu6, Cduiu6, Jduiu6;
wire Qduiu6, Xduiu6, Eeuiu6, Leuiu6, Seuiu6, Zeuiu6, Gfuiu6, Nfuiu6, Ufuiu6, Bguiu6;
wire Iguiu6, Pguiu6, Wguiu6, Dhuiu6, Khuiu6, Rhuiu6, Yhuiu6, Fiuiu6, Miuiu6, Tiuiu6;
wire Ajuiu6, Hjuiu6, Ojuiu6, Vjuiu6, Ckuiu6, Jkuiu6, Qkuiu6, Xkuiu6, Eluiu6, Lluiu6;
wire Sluiu6, Zluiu6, Gmuiu6, Nmuiu6, Umuiu6, Bnuiu6, Inuiu6, Pnuiu6, Wnuiu6, Douiu6;
wire Kouiu6, Rouiu6, Youiu6, Fpuiu6, Mpuiu6, Tpuiu6, Aquiu6, Hquiu6, Oquiu6, Vquiu6;
wire Cruiu6, Jruiu6, Qruiu6, Xruiu6, Esuiu6, Lsuiu6, Ssuiu6, Zsuiu6, Gtuiu6, Ntuiu6;
wire Utuiu6, Buuiu6, Iuuiu6, Puuiu6, Wuuiu6, Dvuiu6, Kvuiu6, Rvuiu6, Yvuiu6, Fwuiu6;
wire Mwuiu6, Twuiu6, Axuiu6, Hxuiu6, Oxuiu6, Vxuiu6, Cyuiu6, Jyuiu6, Qyuiu6, Xyuiu6;
wire Ezuiu6, Lzuiu6, Szuiu6, Zzuiu6, G0viu6, N0viu6, U0viu6, B1viu6, I1viu6, P1viu6;
wire W1viu6, D2viu6, K2viu6, R2viu6, Y2viu6, F3viu6, M3viu6, T3viu6, A4viu6, H4viu6;
wire O4viu6, V4viu6, C5viu6, J5viu6, Q5viu6, X5viu6, E6viu6, L6viu6, S6viu6, Z6viu6;
wire G7viu6, N7viu6, U7viu6, B8viu6, I8viu6, P8viu6, W8viu6, D9viu6, K9viu6, R9viu6;
wire Y9viu6, Faviu6, Maviu6, Taviu6, Abviu6, Hbviu6, Obviu6, Vbviu6, Ccviu6, Jcviu6;
wire Qcviu6, Xcviu6, Edviu6, Ldviu6, Sdviu6, Zdviu6, Geviu6, Neviu6, Ueviu6, Bfviu6;
wire Ifviu6, Pfviu6, Wfviu6, Dgviu6, Kgviu6, Rgviu6, Ygviu6, Fhviu6, Mhviu6, Thviu6;
wire Aiviu6, Hiviu6, Oiviu6, Viviu6, Cjviu6, Jjviu6, Qjviu6, Xjviu6, Ekviu6, Lkviu6;
wire Skviu6, Zkviu6, Glviu6, Nlviu6, Ulviu6, Bmviu6, Imviu6, Pmviu6, Wmviu6, Dnviu6;
wire Knviu6, Rnviu6, Ynviu6, Foviu6, Moviu6, Toviu6, Apviu6, Hpviu6, Opviu6, Vpviu6;
wire Cqviu6, Jqviu6, Qqviu6, Xqviu6, Erviu6, Lrviu6, Srviu6, Zrviu6, Gsviu6, Nsviu6;
wire Usviu6, Btviu6, Itviu6, Ptviu6, Wtviu6, Duviu6, Kuviu6, Ruviu6, Yuviu6, Fvviu6;
wire Mvviu6, Tvviu6, Awviu6, Hwviu6, Owviu6, Vwviu6, Cxviu6, Jxviu6, Qxviu6, Xxviu6;
wire Eyviu6, Lyviu6, Syviu6, Zyviu6, Gzviu6, Nzviu6, Uzviu6, B0wiu6, I0wiu6, P0wiu6;
wire W0wiu6, D1wiu6, K1wiu6, R1wiu6, Y1wiu6, F2wiu6, M2wiu6, T2wiu6, A3wiu6, H3wiu6;
wire O3wiu6, V3wiu6, C4wiu6, J4wiu6, Q4wiu6, X4wiu6, E5wiu6, L5wiu6, S5wiu6, Z5wiu6;
wire G6wiu6, N6wiu6, U6wiu6, B7wiu6, I7wiu6, P7wiu6, W7wiu6, D8wiu6, K8wiu6, R8wiu6;
wire Y8wiu6, F9wiu6, M9wiu6, T9wiu6, Aawiu6, Hawiu6, Oawiu6, Vawiu6, Cbwiu6, Jbwiu6;
wire Qbwiu6, Xbwiu6, Ecwiu6, Lcwiu6, Scwiu6, Zcwiu6, Gdwiu6, Ndwiu6, Udwiu6, Bewiu6;
wire Iewiu6, Pewiu6, Wewiu6, Dfwiu6, Kfwiu6, Rfwiu6, Yfwiu6, Fgwiu6, Mgwiu6, Tgwiu6;
wire Ahwiu6, Hhwiu6, Ohwiu6, Vhwiu6, Ciwiu6, Jiwiu6, Qiwiu6, Xiwiu6, Ejwiu6, Ljwiu6;
wire Sjwiu6, Zjwiu6, Gkwiu6, Nkwiu6, Ukwiu6, Blwiu6, Ilwiu6, Plwiu6, Wlwiu6, Dmwiu6;
wire Kmwiu6, Rmwiu6, Ymwiu6, Fnwiu6, Mnwiu6, Tnwiu6, Aowiu6, Howiu6, Oowiu6, Vowiu6;
wire Cpwiu6, Jpwiu6, Qpwiu6, Xpwiu6, Eqwiu6, Lqwiu6, Sqwiu6, Zqwiu6, Grwiu6, Nrwiu6;
wire Urwiu6, Bswiu6, Iswiu6, Pswiu6, Wswiu6, Dtwiu6, Ktwiu6, Rtwiu6, Ytwiu6, Fuwiu6;
wire Muwiu6, Tuwiu6, Avwiu6, Hvwiu6, Ovwiu6, Vvwiu6, Cwwiu6, Jwwiu6, Qwwiu6, Xwwiu6;
wire Exwiu6, Lxwiu6, Sxwiu6, Zxwiu6, Gywiu6, Nywiu6, Uywiu6, Bzwiu6, Izwiu6, Pzwiu6;
wire Wzwiu6, D0xiu6, K0xiu6, R0xiu6, Y0xiu6, F1xiu6, M1xiu6, T1xiu6, A2xiu6, H2xiu6;
wire O2xiu6, V2xiu6, C3xiu6, J3xiu6, Q3xiu6, X3xiu6, E4xiu6, L4xiu6, S4xiu6, Z4xiu6;
wire G5xiu6, N5xiu6, U5xiu6, B6xiu6, I6xiu6, P6xiu6, W6xiu6, D7xiu6, K7xiu6, R7xiu6;
wire Y7xiu6, F8xiu6, M8xiu6, T8xiu6, A9xiu6, H9xiu6, O9xiu6, V9xiu6, Caxiu6, Jaxiu6;
wire Qaxiu6, Xaxiu6, Ebxiu6, Lbxiu6, Sbxiu6, Zbxiu6, Gcxiu6, Ncxiu6, Ucxiu6, Bdxiu6;
wire Idxiu6, Pdxiu6, Wdxiu6, Dexiu6, Kexiu6, Rexiu6, Yexiu6, Ffxiu6, Mfxiu6, Tfxiu6;
wire Agxiu6, Hgxiu6, Ogxiu6, Vgxiu6, Chxiu6, Jhxiu6, Qhxiu6, Xhxiu6, Eixiu6, Lixiu6;
wire Sixiu6, Zixiu6, Gjxiu6, Njxiu6, Ujxiu6, Bkxiu6, Ikxiu6, Pkxiu6, Wkxiu6, Dlxiu6;
wire Klxiu6, Rlxiu6, Ylxiu6, Fmxiu6, Mmxiu6, Tmxiu6, Anxiu6, Hnxiu6, Onxiu6, Vnxiu6;
wire Coxiu6, Joxiu6, Qoxiu6, Xoxiu6, Epxiu6, Lpxiu6, Spxiu6, Zpxiu6, Gqxiu6, Nqxiu6;
wire Uqxiu6, Brxiu6, Irxiu6, Prxiu6, Wrxiu6, Dsxiu6, Ksxiu6, Rsxiu6, Ysxiu6, Ftxiu6;
wire Mtxiu6, Ttxiu6, Auxiu6, Huxiu6, Ouxiu6, Vuxiu6, Cvxiu6, Jvxiu6, Qvxiu6, Xvxiu6;
wire Ewxiu6, Lwxiu6, Swxiu6, Zwxiu6, Gxxiu6, Nxxiu6, Uxxiu6, Byxiu6, Iyxiu6, Pyxiu6;
wire Wyxiu6, Dzxiu6, Kzxiu6, Rzxiu6, Yzxiu6, F0yiu6, M0yiu6, T0yiu6, A1yiu6, H1yiu6;
wire O1yiu6, V1yiu6, C2yiu6, J2yiu6, Q2yiu6, X2yiu6, E3yiu6, L3yiu6, S3yiu6, Z3yiu6;
wire G4yiu6, N4yiu6, U4yiu6, B5yiu6, I5yiu6, P5yiu6, W5yiu6, D6yiu6, K6yiu6, R6yiu6;
wire Y6yiu6, F7yiu6, M7yiu6, T7yiu6, A8yiu6, H8yiu6, O8yiu6, V8yiu6, C9yiu6, J9yiu6;
wire Q9yiu6, X9yiu6, Eayiu6, Layiu6, Sayiu6, Zayiu6, Gbyiu6, Nbyiu6, Ubyiu6, Bcyiu6;
wire Icyiu6, Pcyiu6, Wcyiu6, Ddyiu6, Kdyiu6, Rdyiu6, Ydyiu6, Feyiu6, Meyiu6, Teyiu6;
wire Afyiu6, Hfyiu6, Ofyiu6, Vfyiu6, Cgyiu6, Jgyiu6, Qgyiu6, Xgyiu6, Ehyiu6, Lhyiu6;
wire Shyiu6, Zhyiu6, Giyiu6, Niyiu6, Uiyiu6, Bjyiu6, Ijyiu6, Pjyiu6, Wjyiu6, Dkyiu6;
wire Kkyiu6, Rkyiu6, Ykyiu6, Flyiu6, Mlyiu6, Tlyiu6, Amyiu6, Hmyiu6, Omyiu6, Vmyiu6;
wire Cnyiu6, Jnyiu6, Qnyiu6, Xnyiu6, Eoyiu6, Loyiu6, Soyiu6, Zoyiu6, Gpyiu6, Npyiu6;
wire Upyiu6, Bqyiu6, Iqyiu6, Pqyiu6, Wqyiu6, Dryiu6, Kryiu6, Rryiu6, Yryiu6, Fsyiu6;
wire Msyiu6, Tsyiu6, Atyiu6, Htyiu6, Otyiu6, Vtyiu6, Cuyiu6, Juyiu6, Quyiu6, Xuyiu6;
wire Evyiu6, Lvyiu6, Svyiu6, Zvyiu6, Gwyiu6, Nwyiu6, Uwyiu6, Bxyiu6, Ixyiu6, Pxyiu6;
wire Wxyiu6, Dyyiu6, Kyyiu6, Ryyiu6, Yyyiu6, Fzyiu6, Mzyiu6, Tzyiu6, A0ziu6, H0ziu6;
wire O0ziu6, V0ziu6, C1ziu6, J1ziu6, Q1ziu6, X1ziu6, E2ziu6, L2ziu6, S2ziu6, Z2ziu6;
wire G3ziu6, N3ziu6, U3ziu6, B4ziu6, I4ziu6, P4ziu6, W4ziu6, D5ziu6, K5ziu6, R5ziu6;
wire Y5ziu6, F6ziu6, M6ziu6, T6ziu6, A7ziu6, H7ziu6, O7ziu6, V7ziu6, C8ziu6, J8ziu6;
wire Q8ziu6, X8ziu6, E9ziu6, L9ziu6, S9ziu6, Z9ziu6, Gaziu6, Naziu6, Uaziu6, Bbziu6;
wire Ibziu6, Pbziu6, Wbziu6, Dcziu6, Kcziu6, Rcziu6, Ycziu6, Fdziu6, Mdziu6, Tdziu6;
wire Aeziu6, Heziu6, Oeziu6, Veziu6, Cfziu6, Jfziu6, Qfziu6, Xfziu6, Egziu6, Lgziu6;
wire Sgziu6, Zgziu6, Ghziu6, Nhziu6, Uhziu6, Biziu6, Iiziu6, Piziu6, Wiziu6, Djziu6;
wire Kjziu6, Rjziu6, Yjziu6, Fkziu6, Mkziu6, Tkziu6, Alziu6, Hlziu6, Olziu6, Vlziu6;
wire Cmziu6, Jmziu6, Qmziu6, Xmziu6, Enziu6, Lnziu6, Snziu6, Znziu6, Goziu6, Noziu6;
wire Uoziu6, Bpziu6, Ipziu6, Ppziu6, Wpziu6, Dqziu6, Kqziu6, Rqziu6, Yqziu6, Frziu6;
wire Mrziu6, Trziu6, Asziu6, Hsziu6, Osziu6, Vsziu6, Ctziu6, Jtziu6, Qtziu6, Xtziu6;
wire Euziu6, Luziu6, Suziu6, Zuziu6, Gvziu6, Nvziu6, Uvziu6, Bwziu6, Iwziu6, Pwziu6;
wire Wwziu6, Dxziu6, Kxziu6, Rxziu6, Yxziu6, Fyziu6, Myziu6, Tyziu6, Azziu6, Hzziu6;
wire Ozziu6, Vzziu6, C00ju6, J00ju6, Q00ju6, X00ju6, E10ju6, L10ju6, S10ju6, Z10ju6;
wire G20ju6, N20ju6, U20ju6, B30ju6, I30ju6, P30ju6, W30ju6, D40ju6, K40ju6, R40ju6;
wire Y40ju6, F50ju6, M50ju6, T50ju6, A60ju6, H60ju6, O60ju6, V60ju6, C70ju6, J70ju6;
wire Q70ju6, X70ju6, E80ju6, L80ju6, S80ju6, Z80ju6, G90ju6, N90ju6, U90ju6, Ba0ju6;
wire Ia0ju6, Pa0ju6, Wa0ju6, Db0ju6, Kb0ju6, Rb0ju6, Yb0ju6, Fc0ju6, Mc0ju6, Tc0ju6;
wire Ad0ju6, Hd0ju6, Od0ju6, Vd0ju6, Ce0ju6, Je0ju6, Qe0ju6, Xe0ju6, Ef0ju6, Lf0ju6;
wire Sf0ju6, Zf0ju6, Gg0ju6, Ng0ju6, Ug0ju6, Bh0ju6, Ih0ju6, Ph0ju6, Wh0ju6, Di0ju6;
wire Ki0ju6, Ri0ju6, Yi0ju6, Fj0ju6, Mj0ju6, Tj0ju6, Ak0ju6, Hk0ju6, Ok0ju6, Vk0ju6;
wire Cl0ju6, Jl0ju6, Ql0ju6, Xl0ju6, Em0ju6, Lm0ju6, Sm0ju6, Zm0ju6, Gn0ju6, Nn0ju6;
wire Un0ju6, Bo0ju6, Io0ju6, Po0ju6, Wo0ju6, Dp0ju6, Kp0ju6, Rp0ju6, Yp0ju6, Fq0ju6;
wire Mq0ju6, Tq0ju6, Ar0ju6, Hr0ju6, Or0ju6, Vr0ju6, Cs0ju6, Js0ju6, Qs0ju6, Xs0ju6;
wire Et0ju6, Lt0ju6, St0ju6, Zt0ju6, Gu0ju6, Nu0ju6, Uu0ju6, Bv0ju6, Iv0ju6, Pv0ju6;
wire Wv0ju6, Dw0ju6, Kw0ju6, Rw0ju6, Yw0ju6, Fx0ju6, Mx0ju6, Tx0ju6, Ay0ju6, Hy0ju6;
wire Oy0ju6, Vy0ju6, Cz0ju6, Jz0ju6, Qz0ju6, Xz0ju6, E01ju6, L01ju6, S01ju6, Z01ju6;
wire G11ju6, N11ju6, U11ju6, B21ju6, I21ju6, P21ju6, W21ju6, D31ju6, K31ju6, R31ju6;
wire Y31ju6, F41ju6, M41ju6, T41ju6, A51ju6, H51ju6, O51ju6, V51ju6, C61ju6, J61ju6;
wire Q61ju6, X61ju6, E71ju6, L71ju6, S71ju6, Z71ju6, G81ju6, N81ju6, U81ju6, B91ju6;
wire I91ju6, P91ju6, W91ju6, Da1ju6, Ka1ju6, Ra1ju6, Ya1ju6, Fb1ju6, Mb1ju6, Tb1ju6;
wire Ac1ju6, Hc1ju6, Oc1ju6, Vc1ju6, Cd1ju6, Jd1ju6, Qd1ju6, Xd1ju6, Ee1ju6, Le1ju6;
wire Se1ju6, Ze1ju6, Gf1ju6, Nf1ju6, Uf1ju6, Bg1ju6, Ig1ju6, Pg1ju6, Wg1ju6, Dh1ju6;
wire Kh1ju6, Rh1ju6, Yh1ju6, Fi1ju6, Mi1ju6, Ti1ju6, Aj1ju6, Hj1ju6, Oj1ju6, Vj1ju6;
wire Ck1ju6, Jk1ju6, Qk1ju6, Xk1ju6, El1ju6, Ll1ju6, Sl1ju6, Zl1ju6, Gm1ju6, Nm1ju6;
wire Um1ju6, Bn1ju6, In1ju6, Pn1ju6, Wn1ju6, Do1ju6, Ko1ju6, Ro1ju6, Yo1ju6, Fp1ju6;
wire Mp1ju6, Tp1ju6, Aq1ju6, Hq1ju6, Oq1ju6, Vq1ju6, Cr1ju6, Jr1ju6, Qr1ju6, Xr1ju6;
wire Es1ju6, Ls1ju6, Ss1ju6, Zs1ju6, Gt1ju6, Nt1ju6, Ut1ju6, Bu1ju6, Iu1ju6, Pu1ju6;
wire Wu1ju6, Dv1ju6, Kv1ju6, Rv1ju6, Yv1ju6, Fw1ju6, Mw1ju6, Tw1ju6, Ax1ju6, Hx1ju6;
wire Ox1ju6, Vx1ju6, Cy1ju6, Jy1ju6, Qy1ju6, Xy1ju6, Ez1ju6, Lz1ju6, Sz1ju6, Zz1ju6;
wire G02ju6, N02ju6, U02ju6, B12ju6, I12ju6, P12ju6, W12ju6, D22ju6, K22ju6, R22ju6;
wire Y22ju6, F32ju6, M32ju6, T32ju6, A42ju6, H42ju6, O42ju6, V42ju6, C52ju6, J52ju6;
wire Q52ju6, X52ju6, E62ju6, L62ju6, S62ju6, Z62ju6, G72ju6, N72ju6, U72ju6, B82ju6;
wire I82ju6, P82ju6, W82ju6, D92ju6, K92ju6, R92ju6, Y92ju6, Fa2ju6, Ma2ju6, Ta2ju6;
wire Ab2ju6, Hb2ju6, Ob2ju6, Vb2ju6, Cc2ju6, Jc2ju6, Qc2ju6, Xc2ju6, Ed2ju6, Ld2ju6;
wire Sd2ju6, Zd2ju6, Ge2ju6, Ne2ju6, Ue2ju6, Bf2ju6, If2ju6, Pf2ju6, Wf2ju6, Dg2ju6;
wire Kg2ju6, Rg2ju6, Yg2ju6, Fh2ju6, Mh2ju6, Th2ju6, Ai2ju6, Hi2ju6, Oi2ju6, Vi2ju6;
wire Cj2ju6, Jj2ju6, Qj2ju6, Xj2ju6, Ek2ju6, Lk2ju6, Sk2ju6, Zk2ju6, Gl2ju6, Nl2ju6;
wire Ul2ju6, Bm2ju6, Im2ju6, Pm2ju6, Wm2ju6, Dn2ju6, Kn2ju6, Rn2ju6, Yn2ju6, Fo2ju6;
wire Mo2ju6, To2ju6, Ap2ju6, Hp2ju6, Op2ju6, Vp2ju6, Cq2ju6, Jq2ju6, Qq2ju6, Xq2ju6;
wire Er2ju6, Lr2ju6, Sr2ju6, Zr2ju6, Gs2ju6, Ns2ju6, Us2ju6, Bt2ju6, It2ju6, Pt2ju6;
wire Wt2ju6, Du2ju6, Ku2ju6, Ru2ju6, Yu2ju6, Fv2ju6, Mv2ju6, Tv2ju6, Aw2ju6, Hw2ju6;
wire Ow2ju6, Vw2ju6, Cx2ju6, Jx2ju6, Qx2ju6, Xx2ju6, Ey2ju6, Ly2ju6, Sy2ju6, Zy2ju6;
wire Gz2ju6, Nz2ju6, Uz2ju6, B03ju6, I03ju6, P03ju6, W03ju6, D13ju6, K13ju6, R13ju6;
wire Y13ju6, F23ju6, M23ju6, T23ju6, A33ju6, H33ju6, O33ju6, V33ju6, C43ju6, J43ju6;
wire Q43ju6, X43ju6, E53ju6, L53ju6, S53ju6, Z53ju6, G63ju6, N63ju6, U63ju6, B73ju6;
wire I73ju6, P73ju6, W73ju6, D83ju6, K83ju6, R83ju6, Y83ju6, F93ju6, M93ju6, T93ju6;
wire Aa3ju6, Ha3ju6, Oa3ju6, Va3ju6, Cb3ju6, Jb3ju6, Qb3ju6, Xb3ju6, Ec3ju6, Lc3ju6;
wire Sc3ju6, Zc3ju6, Gd3ju6, Nd3ju6, Ud3ju6, Be3ju6, Ie3ju6, Pe3ju6, We3ju6, Df3ju6;
wire Kf3ju6, Rf3ju6, Yf3ju6, Fg3ju6, Mg3ju6, Tg3ju6, Ah3ju6, Hh3ju6, Oh3ju6, Vh3ju6;
wire Ci3ju6, Ji3ju6, Qi3ju6, Xi3ju6, Ej3ju6, Lj3ju6, Sj3ju6, Zj3ju6, Gk3ju6, Nk3ju6;
wire Uk3ju6, Bl3ju6, Il3ju6, Pl3ju6, Wl3ju6, Dm3ju6, Km3ju6, Rm3ju6, Ym3ju6, Fn3ju6;
wire Mn3ju6, Tn3ju6, Ao3ju6, Ho3ju6, Oo3ju6, Vo3ju6, Cp3ju6, Jp3ju6, Qp3ju6, Xp3ju6;
wire Eq3ju6, Lq3ju6, Sq3ju6, Zq3ju6, Gr3ju6, Nr3ju6, Ur3ju6, Bs3ju6, Is3ju6, Ps3ju6;
wire Ws3ju6, Dt3ju6, Kt3ju6, Rt3ju6, Yt3ju6, Fu3ju6, Mu3ju6, Tu3ju6, Av3ju6, Hv3ju6;
wire Ov3ju6, Vv3ju6, Cw3ju6, Jw3ju6, Qw3ju6, Xw3ju6, Ex3ju6, Lx3ju6, Sx3ju6, Zx3ju6;
wire Gy3ju6, Ny3ju6, Uy3ju6, Bz3ju6, Iz3ju6, Pz3ju6, Wz3ju6, D04ju6, K04ju6, R04ju6;
wire Y04ju6, F14ju6, M14ju6, T14ju6, A24ju6, H24ju6, O24ju6, V24ju6, C34ju6, J34ju6;
wire Q34ju6, X34ju6, E44ju6, L44ju6, S44ju6, Z44ju6, G54ju6, N54ju6, U54ju6, B64ju6;
wire I64ju6, P64ju6, W64ju6, D74ju6, K74ju6, R74ju6, Y74ju6, F84ju6, M84ju6, T84ju6;
wire A94ju6, H94ju6, O94ju6, V94ju6, Ca4ju6, Ja4ju6, Qa4ju6, Xa4ju6, Eb4ju6, Lb4ju6;
wire Sb4ju6, Zb4ju6, Gc4ju6, Nc4ju6, Uc4ju6, Bd4ju6, Id4ju6, Pd4ju6, Wd4ju6, De4ju6;
wire Ke4ju6, Re4ju6, Ye4ju6, Ff4ju6, Mf4ju6, Tf4ju6, Ag4ju6, Hg4ju6, Og4ju6, Vg4ju6;
wire Ch4ju6, Jh4ju6, Qh4ju6, Xh4ju6, Ei4ju6, Li4ju6, Si4ju6, Zi4ju6, Gj4ju6, Nj4ju6;
wire Uj4ju6, Bk4ju6, Ik4ju6, Pk4ju6, Wk4ju6, Dl4ju6, Kl4ju6, Rl4ju6, Yl4ju6, Fm4ju6;
wire Mm4ju6, Tm4ju6, An4ju6, Hn4ju6, On4ju6, Vn4ju6, Co4ju6, Jo4ju6, Qo4ju6, Xo4ju6;
wire Ep4ju6, Lp4ju6, Sp4ju6, Zp4ju6, Gq4ju6, Nq4ju6, Uq4ju6, Br4ju6, Ir4ju6, Pr4ju6;
wire Wr4ju6, Ds4ju6, Ks4ju6, Rs4ju6, Ys4ju6, Ft4ju6, Mt4ju6, Tt4ju6, Au4ju6, Hu4ju6;
wire Ou4ju6, Vu4ju6, Cv4ju6, Jv4ju6, Qv4ju6, Xv4ju6, Ew4ju6, Lw4ju6, Sw4ju6, Zw4ju6;
wire Gx4ju6, Nx4ju6, Ux4ju6, By4ju6, Iy4ju6, Py4ju6, Wy4ju6, Dz4ju6, Kz4ju6, Rz4ju6;
wire Yz4ju6, F05ju6, M05ju6, T05ju6, A15ju6, H15ju6, O15ju6, V15ju6, C25ju6, J25ju6;
wire Q25ju6, X25ju6, E35ju6, L35ju6, S35ju6, Z35ju6, G45ju6, N45ju6, U45ju6, B55ju6;
wire I55ju6, P55ju6, W55ju6, D65ju6, K65ju6, R65ju6, Y65ju6, F75ju6, M75ju6, T75ju6;
wire A85ju6, H85ju6, O85ju6, V85ju6, C95ju6, J95ju6, Q95ju6, X95ju6, Ea5ju6, La5ju6;
wire Sa5ju6, Za5ju6, Gb5ju6, Nb5ju6, Ub5ju6, Bc5ju6, Ic5ju6, Pc5ju6, Wc5ju6, Dd5ju6;
wire Kd5ju6, Rd5ju6, Yd5ju6, Fe5ju6, Me5ju6, Te5ju6, Af5ju6, Hf5ju6, Of5ju6, Vf5ju6;
wire Cg5ju6, Jg5ju6, Qg5ju6, Xg5ju6, Eh5ju6, Lh5ju6, Sh5ju6, Zh5ju6, Gi5ju6, Ni5ju6;
wire Ui5ju6, Bj5ju6, Ij5ju6, Pj5ju6, Wj5ju6, Dk5ju6, Kk5ju6, Rk5ju6, Yk5ju6, Fl5ju6;
wire Ml5ju6, Tl5ju6, Am5ju6, Hm5ju6, Om5ju6, Vm5ju6, Cn5ju6, Jn5ju6, Qn5ju6, Xn5ju6;
wire Eo5ju6, Lo5ju6, So5ju6, Zo5ju6, Gp5ju6, Np5ju6, Up5ju6, Bq5ju6, Iq5ju6, Pq5ju6;
wire Wq5ju6, Dr5ju6, Kr5ju6, Rr5ju6, Yr5ju6, Fs5ju6, Ms5ju6, Ts5ju6, At5ju6, Ht5ju6;
wire Ot5ju6, Vt5ju6, Cu5ju6, Ju5ju6, Qu5ju6, Xu5ju6, Ev5ju6, Lv5ju6, Sv5ju6, Zv5ju6;
wire Gw5ju6, Nw5ju6, Uw5ju6, Bx5ju6, Ix5ju6, Px5ju6, Wx5ju6, Dy5ju6, Ky5ju6, Ry5ju6;
wire Yy5ju6, Fz5ju6, Mz5ju6, Tz5ju6, A06ju6, H06ju6, O06ju6, V06ju6, C16ju6, J16ju6;
wire Q16ju6, X16ju6, E26ju6, L26ju6, S26ju6, Z26ju6, G36ju6, N36ju6, U36ju6, B46ju6;
wire I46ju6, P46ju6, W46ju6, D56ju6, K56ju6, R56ju6, Y56ju6, F66ju6, M66ju6, T66ju6;
wire A76ju6, H76ju6, O76ju6, V76ju6, C86ju6, J86ju6, Q86ju6, X86ju6, E96ju6, L96ju6;
wire S96ju6, Z96ju6, Ga6ju6, Na6ju6, Ua6ju6, Bb6ju6, Ib6ju6, Pb6ju6, Wb6ju6, Dc6ju6;
wire Kc6ju6, Rc6ju6, Yc6ju6, Fd6ju6, Md6ju6, Td6ju6, Ae6ju6, He6ju6, Oe6ju6, Ve6ju6;
wire Cf6ju6, Jf6ju6, Qf6ju6, Xf6ju6, Eg6ju6, Lg6ju6, Sg6ju6, Zg6ju6, Gh6ju6, Nh6ju6;
wire Uh6ju6, Bi6ju6, Ii6ju6, Pi6ju6, Wi6ju6, Dj6ju6, Kj6ju6, Rj6ju6, Yj6ju6, Fk6ju6;
wire Mk6ju6, Tk6ju6, Al6ju6, Hl6ju6, Ol6ju6, Vl6ju6, Cm6ju6, Jm6ju6, Qm6ju6, Xm6ju6;
wire En6ju6, Ln6ju6, Sn6ju6, Zn6ju6, Go6ju6, No6ju6, Uo6ju6, Bp6ju6, Ip6ju6, Pp6ju6;
wire Wp6ju6, Dq6ju6, Kq6ju6, Rq6ju6, Yq6ju6, Fr6ju6, Mr6ju6, Tr6ju6, As6ju6, Hs6ju6;
wire Os6ju6, Vs6ju6, Ct6ju6, Jt6ju6, Qt6ju6, Xt6ju6, Eu6ju6, Lu6ju6, Su6ju6, Zu6ju6;
wire Gv6ju6, Nv6ju6, Uv6ju6, Bw6ju6, Iw6ju6, Pw6ju6, Ww6ju6, Dx6ju6, Kx6ju6, Rx6ju6;
wire Yx6ju6, Fy6ju6, My6ju6, Ty6ju6, Az6ju6, Hz6ju6, Oz6ju6, Vz6ju6, C07ju6, J07ju6;
wire Q07ju6, X07ju6, E17ju6, L17ju6, S17ju6, Z17ju6, G27ju6, N27ju6, U27ju6, B37ju6;
wire I37ju6, P37ju6, W37ju6, D47ju6, K47ju6, R47ju6, Y47ju6, F57ju6, M57ju6, T57ju6;
wire A67ju6, H67ju6, O67ju6, V67ju6, C77ju6, J77ju6, Q77ju6, X77ju6, E87ju6, L87ju6;
wire S87ju6, Z87ju6, G97ju6, N97ju6, U97ju6, Ba7ju6, Ia7ju6, Pa7ju6, Wa7ju6, Db7ju6;
wire Kb7ju6, Rb7ju6, Yb7ju6, Fc7ju6, Mc7ju6, Tc7ju6, Ad7ju6, Hd7ju6, Od7ju6, Vd7ju6;
wire Ce7ju6, Je7ju6, Qe7ju6, Xe7ju6, Ef7ju6, Lf7ju6, Sf7ju6, Zf7ju6, Gg7ju6, Ng7ju6;
wire Ug7ju6, Bh7ju6, Ih7ju6, Ph7ju6, Wh7ju6, Di7ju6, Ki7ju6, Ri7ju6, Yi7ju6, Fj7ju6;
wire Mj7ju6, Tj7ju6, Ak7ju6, Hk7ju6, Ok7ju6, Vk7ju6, Cl7ju6, Jl7ju6, Ql7ju6, Xl7ju6;
wire Em7ju6, Lm7ju6, Sm7ju6, Zm7ju6, Gn7ju6, Nn7ju6, Un7ju6, Bo7ju6, Io7ju6, Po7ju6;
wire Wo7ju6, Dp7ju6, Kp7ju6, Rp7ju6, Yp7ju6, Fq7ju6, Mq7ju6, Tq7ju6, Ar7ju6, Hr7ju6;
wire Or7ju6, Vr7ju6, Cs7ju6, Js7ju6, Qs7ju6, Xs7ju6, Et7ju6, Lt7ju6, St7ju6, Zt7ju6;
wire Gu7ju6, Nu7ju6, Uu7ju6, Bv7ju6, Iv7ju6, Pv7ju6, Wv7ju6, Dw7ju6, Kw7ju6, Rw7ju6;
wire Yw7ju6, Fx7ju6, Mx7ju6, Tx7ju6, Ay7ju6, Hy7ju6, Oy7ju6, Vy7ju6, Cz7ju6, Jz7ju6;
wire Qz7ju6, Xz7ju6, E08ju6, L08ju6, S08ju6, Z08ju6, G18ju6, N18ju6, U18ju6, B28ju6;
wire I28ju6, P28ju6, W28ju6, D38ju6, K38ju6, R38ju6, Y38ju6, F48ju6, M48ju6, T48ju6;
wire A58ju6, H58ju6, O58ju6, V58ju6, C68ju6, J68ju6, Q68ju6, X68ju6, E78ju6, L78ju6;
wire S78ju6, Z78ju6, G88ju6, N88ju6, U88ju6, B98ju6, I98ju6, P98ju6, W98ju6, Da8ju6;
wire Ka8ju6, Ra8ju6, Ya8ju6, Fb8ju6, Mb8ju6, Tb8ju6, Ac8ju6, Hc8ju6, Oc8ju6, Vc8ju6;
wire Cd8ju6, Jd8ju6, Qd8ju6, Xd8ju6, Ee8ju6, Le8ju6, Se8ju6, Ze8ju6, Gf8ju6, Nf8ju6;
wire Uf8ju6, Bg8ju6, Ig8ju6, Pg8ju6, Wg8ju6, Dh8ju6, Kh8ju6, Rh8ju6, Yh8ju6, Fi8ju6;
wire Mi8ju6, Ti8ju6, Aj8ju6, Hj8ju6, Oj8ju6, Vj8ju6, Ck8ju6, Jk8ju6, Qk8ju6, Xk8ju6;
wire El8ju6, Ll8ju6, Sl8ju6, Zl8ju6, Gm8ju6, Nm8ju6, Um8ju6, Bn8ju6, In8ju6, Pn8ju6;
wire Wn8ju6, Do8ju6, Ko8ju6, Ro8ju6, Yo8ju6, Fp8ju6, Mp8ju6, Tp8ju6, Aq8ju6, Hq8ju6;
wire Oq8ju6, Vq8ju6, Cr8ju6, Jr8ju6, Qr8ju6, Xr8ju6, Es8ju6, Ls8ju6, Ss8ju6, Zs8ju6;
wire Gt8ju6, Nt8ju6, Ut8ju6, Bu8ju6, Iu8ju6, Pu8ju6, Wu8ju6, Dv8ju6, Kv8ju6, Rv8ju6;
wire Yv8ju6, Fw8ju6, Mw8ju6, Tw8ju6, Ax8ju6, Hx8ju6, Ox8ju6, Vx8ju6, Cy8ju6, Jy8ju6;
wire Qy8ju6, Xy8ju6, Ez8ju6, Lz8ju6, Sz8ju6, Zz8ju6, G09ju6, N09ju6, U09ju6, B19ju6;
wire I19ju6, P19ju6, W19ju6, D29ju6, K29ju6, R29ju6, Y29ju6, F39ju6, M39ju6, T39ju6;
wire A49ju6, H49ju6, O49ju6, V49ju6, C59ju6, J59ju6, Q59ju6, X59ju6, E69ju6, L69ju6;
wire S69ju6, Z69ju6, G79ju6, N79ju6, U79ju6, B89ju6, I89ju6, P89ju6, W89ju6, D99ju6;
wire K99ju6, R99ju6, Y99ju6, Fa9ju6, Ma9ju6, Ta9ju6, Ab9ju6, Hb9ju6, Ob9ju6, Vb9ju6;
wire Cc9ju6, Jc9ju6, Qc9ju6, Xc9ju6, Ed9ju6, Ld9ju6, Sd9ju6, Zd9ju6, Ge9ju6, Ne9ju6;
wire Ue9ju6, Bf9ju6, If9ju6, Pf9ju6, Wf9ju6, Dg9ju6, Kg9ju6, Rg9ju6, Yg9ju6, Fh9ju6;
wire Mh9ju6, Th9ju6, Ai9ju6, Hi9ju6, Oi9ju6, Vi9ju6, Cj9ju6, Jj9ju6, Qj9ju6, Xj9ju6;
wire Ek9ju6, Lk9ju6, Sk9ju6, Zk9ju6, Gl9ju6, Nl9ju6, Ul9ju6, Bm9ju6, Im9ju6, Pm9ju6;
wire Wm9ju6, Dn9ju6, Kn9ju6, Rn9ju6, Yn9ju6, Fo9ju6, Mo9ju6, To9ju6, Ap9ju6, Hp9ju6;
wire Op9ju6, Vp9ju6, Cq9ju6, Jq9ju6, Qq9ju6, Xq9ju6, Er9ju6, Lr9ju6, Sr9ju6, Zr9ju6;
wire Gs9ju6, Ns9ju6, Us9ju6, Bt9ju6, It9ju6, Pt9ju6, Wt9ju6, Du9ju6, Ku9ju6, Ru9ju6;
wire Yu9ju6, Fv9ju6, Mv9ju6, Tv9ju6, Aw9ju6, Hw9ju6, Ow9ju6, Vw9ju6, Cx9ju6, Jx9ju6;
wire Qx9ju6, Xx9ju6, Ey9ju6, Ly9ju6, Sy9ju6, Zy9ju6, Gz9ju6, Nz9ju6, Uz9ju6, B0aju6;
wire I0aju6, P0aju6, W0aju6, D1aju6, K1aju6, R1aju6, Y1aju6, F2aju6, M2aju6, T2aju6;
wire A3aju6, H3aju6, O3aju6, V3aju6, C4aju6, J4aju6, Q4aju6, X4aju6, E5aju6, L5aju6;
wire S5aju6, Z5aju6, G6aju6, N6aju6, U6aju6, B7aju6, I7aju6, P7aju6, W7aju6, D8aju6;
wire K8aju6, R8aju6, Y8aju6, F9aju6, M9aju6, T9aju6, Aaaju6, Haaju6, Oaaju6, Vaaju6;
wire Cbaju6, Jbaju6, Qbaju6, Xbaju6, Ecaju6, Lcaju6, Scaju6, Zcaju6, Gdaju6, Ndaju6;
wire Udaju6, Beaju6, Ieaju6, Peaju6, Weaju6, Dfaju6, Kfaju6, Rfaju6, Yfaju6, Fgaju6;
wire Mgaju6, Tgaju6, Ahaju6, Hhaju6, Ohaju6, Vhaju6, Ciaju6, Jiaju6, Qiaju6, Xiaju6;
wire Ejaju6, Ljaju6, Sjaju6, Zjaju6, Gkaju6, Nkaju6, Ukaju6, Blaju6, Ilaju6, Plaju6;
wire Wlaju6, Dmaju6, Kmaju6, Rmaju6, Ymaju6, Fnaju6, Mnaju6, Tnaju6, Aoaju6, Hoaju6;
wire Ooaju6, Voaju6, Cpaju6, Jpaju6, Qpaju6, Xpaju6, Eqaju6, Lqaju6, Sqaju6, Zqaju6;
wire Graju6, Nraju6, Uraju6, Bsaju6, Isaju6, Psaju6, Wsaju6, Dtaju6, K76ow6, R76ow6;
wire Y76ow6, F86ow6, M86ow6, T86ow6, A96ow6, H96ow6, O96ow6, V96ow6, Ca6ow6, Ja6ow6;
wire Qa6ow6, Xa6ow6, Eb6ow6, Lb6ow6, Sb6ow6, Zb6ow6, Gc6ow6, Nc6ow6, Uc6ow6, Bd6ow6;
wire Id6ow6, Pd6ow6, Wd6ow6, De6ow6, Ke6ow6, Re6ow6, Ye6ow6, Ff6ow6, Mf6ow6, Tf6ow6;
wire Ag6ow6, Hg6ow6, Og6ow6, Vg6ow6, Ch6ow6, Jh6ow6, Qh6ow6, Xh6ow6, Ei6ow6, Li6ow6;
wire Si6ow6, Zi6ow6, Gj6ow6, Nj6ow6, Uj6ow6, Bk6ow6, Ik6ow6, Pk6ow6, Wk6ow6, Dl6ow6;
wire Kl6ow6, Rl6ow6, Yl6ow6, Fm6ow6, Mm6ow6, Tm6ow6, An6ow6, Hn6ow6, On6ow6, Vn6ow6;
wire Co6ow6, Jo6ow6, Qo6ow6, Xo6ow6, Ep6ow6, Lp6ow6, Sp6ow6, Zp6ow6, Gq6ow6, Nq6ow6;
wire Uq6ow6, Br6ow6, Ir6ow6, Pr6ow6, Wr6ow6, Ds6ow6, Ks6ow6, Rs6ow6, Ys6ow6, Ft6ow6;
wire Mt6ow6, Tt6ow6, Au6ow6, Hu6ow6, Ou6ow6, Vu6ow6, Cv6ow6, Jv6ow6, Qv6ow6, Xv6ow6;
wire Ew6ow6, Lw6ow6, Sw6ow6, Zw6ow6, Gx6ow6, Nx6ow6, Ux6ow6, By6ow6, Iy6ow6, Py6ow6;
wire Wy6ow6, Dz6ow6, Kz6ow6, Rz6ow6, Yz6ow6, F07ow6, M07ow6, T07ow6, A17ow6, H17ow6;
wire O17ow6, V17ow6, C27ow6, J27ow6, Q27ow6, X27ow6, E37ow6, L37ow6, S37ow6, Z37ow6;
wire G47ow6, N47ow6, U47ow6, B57ow6, I57ow6, P57ow6, W57ow6, D67ow6, K67ow6, R67ow6;
wire Y67ow6, F77ow6, M77ow6, T77ow6, A87ow6, H87ow6, O87ow6, V87ow6, C97ow6, J97ow6;
wire Q97ow6, X97ow6, Ea7ow6, La7ow6, Sa7ow6, Za7ow6, Gb7ow6, Nb7ow6, Ub7ow6, Bc7ow6;
wire Ic7ow6, Pc7ow6, Wc7ow6, Dd7ow6, Kd7ow6, Rd7ow6, Yd7ow6, Fe7ow6, Me7ow6, Te7ow6;
wire Af7ow6, Hf7ow6, Of7ow6, Vf7ow6, Cg7ow6, Jg7ow6, Qg7ow6, Xg7ow6, Eh7ow6, Lh7ow6;
wire Sh7ow6, Zh7ow6, Gi7ow6, Ni7ow6, Ui7ow6, Bj7ow6, Ij7ow6, Pj7ow6, Wj7ow6, Dk7ow6;
wire Kk7ow6, Rk7ow6, Yk7ow6, Fl7ow6, Ml7ow6, Tl7ow6, Am7ow6, Hm7ow6, Om7ow6, Vm7ow6;
wire Cn7ow6, Jn7ow6, Qn7ow6, Xn7ow6, Eo7ow6, Lo7ow6, So7ow6, Zo7ow6, Gp7ow6, Np7ow6;
wire Up7ow6, Bq7ow6, Iq7ow6, Pq7ow6, Wq7ow6, Dr7ow6, Kr7ow6, Rr7ow6, Yr7ow6, Fs7ow6;
wire Ms7ow6, Ts7ow6, At7ow6, Ht7ow6, Ot7ow6, Vt7ow6, Cu7ow6, Ju7ow6, Qu7ow6, Xu7ow6;
wire Ev7ow6, Lv7ow6, Sv7ow6, Zv7ow6, Gw7ow6, Nw7ow6, Uw7ow6, Bx7ow6, Ix7ow6, Px7ow6;
wire Wx7ow6, Dy7ow6, Ky7ow6, Ry7ow6, Yy7ow6, Fz7ow6, Mz7ow6, Tz7ow6, A08ow6, H08ow6;
wire O08ow6, V08ow6, C18ow6, J18ow6, Q18ow6, X18ow6, E28ow6, L28ow6, S28ow6, Z28ow6;
wire G38ow6, N38ow6, U38ow6, B48ow6, I48ow6, P48ow6, W48ow6, D58ow6, K58ow6, R58ow6;
wire Y58ow6, F68ow6, M68ow6, T68ow6, A78ow6, H78ow6, O78ow6, V78ow6, C88ow6, J88ow6;
wire Q88ow6, X88ow6, E98ow6, L98ow6, S98ow6, Z98ow6, Ga8ow6, Na8ow6, Ua8ow6, Bb8ow6;
wire Ib8ow6, Pb8ow6, Wb8ow6, Dc8ow6, Kc8ow6, Rc8ow6, Yc8ow6, Fd8ow6, Md8ow6, Td8ow6;
wire Ae8ow6, He8ow6, Oe8ow6, Ve8ow6, Cf8ow6, Jf8ow6, Qf8ow6, Xf8ow6, Eg8ow6, Lg8ow6;
wire Sg8ow6, Zg8ow6, Gh8ow6, Nh8ow6, Uh8ow6, Bi8ow6, Ii8ow6, Pi8ow6, Wi8ow6, Dj8ow6;
wire Kj8ow6, Rj8ow6, Yj8ow6, Fk8ow6, Mk8ow6, Tk8ow6, Al8ow6, Hl8ow6, Ol8ow6, Vl8ow6;
wire Cm8ow6, Jm8ow6, Qm8ow6, Xm8ow6, En8ow6, Ln8ow6, Sn8ow6, Zn8ow6, Go8ow6, No8ow6;
wire Uo8ow6, Bp8ow6, Ip8ow6, Pp8ow6, Wp8ow6, Dq8ow6, Kq8ow6, Rq8ow6, Yq8ow6, Fr8ow6;
wire Mr8ow6, Tr8ow6, As8ow6, Hs8ow6, Os8ow6, Vs8ow6, Ct8ow6, Jt8ow6, Qt8ow6, Xt8ow6;
wire Eu8ow6, Lu8ow6, Su8ow6, Zu8ow6, Gv8ow6, Nv8ow6, Uv8ow6, Bw8ow6, Iw8ow6, Pw8ow6;
wire Ww8ow6, Dx8ow6, Kx8ow6, Rx8ow6, Yx8ow6, Fy8ow6, My8ow6, Ty8ow6, Az8ow6, Hz8ow6;
wire Oz8ow6, Vz8ow6, C09ow6, J09ow6, Q09ow6, X09ow6, E19ow6, L19ow6, S19ow6, Z19ow6;
wire G29ow6, N29ow6, U29ow6, B39ow6, I39ow6, P39ow6, W39ow6, D49ow6, K49ow6, R49ow6;
wire Y49ow6, F59ow6, M59ow6, T59ow6, A69ow6, H69ow6, O69ow6, V69ow6, C79ow6, J79ow6;
wire Q79ow6, X79ow6, E89ow6, L89ow6, S89ow6, Z89ow6, G99ow6, N99ow6, U99ow6, Ba9ow6;
wire Ia9ow6, Pa9ow6, Wa9ow6, Db9ow6, Kb9ow6, Rb9ow6, Yb9ow6, Fc9ow6, Mc9ow6, Tc9ow6;
wire Ad9ow6, Hd9ow6, Od9ow6, Vd9ow6, Ce9ow6, Je9ow6, Qe9ow6, Xe9ow6, Ef9ow6, Lf9ow6;
wire Sf9ow6, Zf9ow6, Gg9ow6, Ng9ow6, Ug9ow6, Bh9ow6, Ih9ow6, Ph9ow6, Wh9ow6, Di9ow6;
wire Ki9ow6, Ri9ow6, Yi9ow6, Fj9ow6, Mj9ow6, Tj9ow6, Ak9ow6, Hk9ow6, Ok9ow6, Vk9ow6;
wire Cl9ow6, Jl9ow6, Ql9ow6, Xl9ow6, Em9ow6, Lm9ow6, Sm9ow6, Zm9ow6, Gn9ow6, Nn9ow6;
wire Un9ow6, Bo9ow6, Io9ow6, Po9ow6, Wo9ow6, Dp9ow6, Kp9ow6, Rp9ow6, Yp9ow6, Fq9ow6;
wire Mq9ow6, Tq9ow6, Ar9ow6, Hr9ow6, Or9ow6, Vr9ow6, Cs9ow6, Js9ow6, Qs9ow6, Xs9ow6;
wire Et9ow6, Lt9ow6, St9ow6, Zt9ow6, Gu9ow6, Nu9ow6, Uu9ow6, Bv9ow6, Iv9ow6, Pv9ow6;
wire Wv9ow6, Dw9ow6, Kw9ow6, Rw9ow6, Yw9ow6, Fx9ow6, Mx9ow6, Tx9ow6, Ay9ow6, Hy9ow6;
wire Oy9ow6, Vy9ow6, Cz9ow6, Jz9ow6, Qz9ow6, Xz9ow6, E0aow6, L0aow6, S0aow6, Z0aow6;
wire G1aow6, N1aow6, U1aow6, B2aow6, I2aow6, P2aow6, W2aow6, D3aow6, K3aow6, R3aow6;
wire Y3aow6, F4aow6, M4aow6, T4aow6, A5aow6, H5aow6, O5aow6, V5aow6, C6aow6, J6aow6;
wire Q6aow6, X6aow6, E7aow6, L7aow6, S7aow6, Z7aow6, G8aow6, N8aow6, U8aow6, B9aow6;
wire I9aow6, P9aow6, W9aow6, Daaow6, Kaaow6, Raaow6, Yaaow6, Fbaow6, Mbaow6, Tbaow6;
wire Acaow6, Hcaow6, Ocaow6, Vcaow6, Cdaow6, Jdaow6, Qdaow6, Xdaow6, Eeaow6, Leaow6;
wire Seaow6, Zeaow6, Gfaow6, Nfaow6, Ufaow6, Bgaow6, Igaow6, Pgaow6, Wgaow6, Dhaow6;
wire Khaow6, Rhaow6, Yhaow6, Fiaow6, Miaow6, Tiaow6, Ajaow6, Hjaow6, Ojaow6, Vjaow6;
wire Ckaow6, Jkaow6, Qkaow6, Xkaow6, Elaow6, Llaow6, Slaow6, Zlaow6, Gmaow6, Nmaow6;
wire Umaow6, Bnaow6, Inaow6, Pnaow6, Wnaow6, Doaow6, Koaow6, Roaow6, Yoaow6, Fpaow6;
wire Mpaow6, Tpaow6, Aqaow6, Hqaow6, Oqaow6, Vqaow6, Craow6, Jraow6, Qraow6, Xraow6;
wire Esaow6, Lsaow6, Ssaow6, Zsaow6, Gtaow6, Ntaow6, Utaow6, Buaow6, Iuaow6, Puaow6;
wire Wuaow6, Dvaow6, Kvaow6, Rvaow6, Yvaow6, Fwaow6, Mwaow6, Twaow6, Axaow6, Hxaow6;
wire Oxaow6, Vxaow6, Cyaow6, Jyaow6, Qyaow6, Xyaow6, Ezaow6, Lzaow6, Szaow6, Zzaow6;
wire G0bow6, N0bow6, U0bow6, B1bow6, I1bow6, P1bow6, W1bow6, D2bow6, K2bow6, R2bow6;
wire Y2bow6, F3bow6, M3bow6, T3bow6, A4bow6, H4bow6, O4bow6, V4bow6, C5bow6, J5bow6;
wire Q5bow6, X5bow6, E6bow6, L6bow6, S6bow6, Z6bow6, G7bow6, N7bow6, U7bow6, B8bow6;
wire I8bow6, P8bow6, W8bow6, D9bow6, K9bow6, R9bow6, Y9bow6, Fabow6, Mabow6, Tabow6;
wire Abbow6, Hbbow6, Obbow6, Vbbow6, Ccbow6, Jcbow6, Qcbow6, Xcbow6, Edbow6, Ldbow6;
wire Sdbow6, Zdbow6, Gebow6, Nebow6, Uebow6, Bfbow6, Ifbow6, Pfbow6, Wfbow6, Dgbow6;
wire Kgbow6, Rgbow6, Ygbow6, Fhbow6, Mhbow6, Thbow6, Aibow6, Hibow6, Oibow6, Vibow6;
wire Cjbow6, Jjbow6, Qjbow6, Xjbow6, Ekbow6, Lkbow6, Skbow6, Zkbow6, Glbow6, Nlbow6;
wire Ulbow6, Bmbow6, Imbow6, Pmbow6, Wmbow6, Dnbow6, Knbow6, Rnbow6, Ynbow6, Fobow6;
wire Mobow6, Tobow6, Apbow6, Hpbow6, Opbow6, Vpbow6, Cqbow6, Jqbow6, Qqbow6, Xqbow6;
wire Erbow6, Lrbow6, Srbow6, Zrbow6, Gsbow6, Nsbow6, Usbow6, Btbow6, Itbow6, Ptbow6;
wire Wtbow6, Dubow6, Kubow6, Rubow6, Yubow6, Fvbow6, Mvbow6, Tvbow6, Awbow6, Hwbow6;
wire Owbow6, Vwbow6, Cxbow6, Jxbow6, Qxbow6, Xxbow6, Eybow6, Lybow6, Sybow6, Zybow6;
wire Gzbow6, Nzbow6, Uzbow6, B0cow6, I0cow6, P0cow6, W0cow6, D1cow6, K1cow6, R1cow6;
wire Y1cow6, F2cow6, M2cow6, T2cow6, A3cow6, H3cow6, O3cow6, V3cow6, C4cow6, J4cow6;
wire Q4cow6, X4cow6, E5cow6, L5cow6, S5cow6, Z5cow6, G6cow6, N6cow6, U6cow6, B7cow6;
wire I7cow6, P7cow6, W7cow6, D8cow6, K8cow6, R8cow6, Y8cow6, F9cow6, M9cow6, T9cow6;
wire Aacow6, Hacow6, Oacow6, Vacow6, Cbcow6, Jbcow6, Qbcow6, Xbcow6, Eccow6, Lccow6;
wire Sccow6, Zccow6, Gdcow6, Ndcow6, Udcow6, Becow6, Iecow6, Pecow6, Wecow6, Dfcow6;
wire Kfcow6, Rfcow6, Yfcow6, Fgcow6, Mgcow6, Tgcow6, Ahcow6, Hhcow6, Ohcow6, Vhcow6;
wire Cicow6, Jicow6, Qicow6, Xicow6, Ejcow6, Ljcow6, Sjcow6, Zjcow6, Gkcow6, Nkcow6;
wire Ukcow6, Blcow6, Ilcow6, Plcow6, Wlcow6, Dmcow6, Kmcow6, Rmcow6, Ymcow6, Fncow6;
wire Mncow6, Tncow6, Aocow6, Hocow6, Oocow6, Vocow6, Cpcow6, Jpcow6, Qpcow6, Xpcow6;
wire Eqcow6, Lqcow6, Sqcow6, Zqcow6, Grcow6, Nrcow6, Urcow6, Bscow6, Iscow6, Pscow6;
wire Wscow6, Dtcow6, Ktcow6, Rtcow6, Ytcow6, Fucow6, Mucow6, Tucow6, Avcow6, Hvcow6;
wire Ovcow6, Vvcow6, Cwcow6, Jwcow6, Qwcow6, Xwcow6, Excow6, Lxcow6, Sxcow6, Zxcow6;
wire Gycow6, Nycow6, Uycow6, Bzcow6, Izcow6, Pzcow6, Wzcow6, D0dow6, K0dow6, R0dow6;
wire Y0dow6, F1dow6, M1dow6, T1dow6, A2dow6, H2dow6, O2dow6, V2dow6, C3dow6, J3dow6;
wire Q3dow6, X3dow6, E4dow6, L4dow6, S4dow6, Z4dow6, G5dow6, N5dow6, U5dow6, B6dow6;
wire I6dow6, P6dow6, W6dow6, D7dow6, K7dow6, R7dow6, Y7dow6, F8dow6, M8dow6, T8dow6;
wire A9dow6, H9dow6, O9dow6, V9dow6, Cadow6, Jadow6, Qadow6, Xadow6, Ebdow6, Lbdow6;
wire Sbdow6, Zbdow6, Gcdow6, Ncdow6, Ucdow6, Bddow6, Iddow6, Pddow6, Wddow6, Dedow6;
wire Kedow6, Redow6, Yedow6, Ffdow6, Mfdow6, Tfdow6, Agdow6, Hgdow6, Ogdow6, Vgdow6;
wire Chdow6, Jhdow6, Qhdow6, Xhdow6, Eidow6, Lidow6, Sidow6, Zidow6, Gjdow6, Njdow6;
wire Ujdow6, Bkdow6, Ikdow6, Pkdow6, Wkdow6, Dldow6, Kldow6, Rldow6, Yldow6, Fmdow6;
wire Mmdow6, Tmdow6, Andow6, Hndow6, Ondow6, Vndow6, Codow6, Jodow6, Qodow6, Xodow6;
wire Epdow6, Lpdow6, Spdow6, Zpdow6, Gqdow6, Nqdow6, Uqdow6, Brdow6, Irdow6, Prdow6;
wire Wrdow6, Dsdow6, Ksdow6, Rsdow6, Ysdow6, Ftdow6, Mtdow6, Ttdow6, Audow6, Hudow6;
wire Oudow6, Vudow6, Cvdow6, Jvdow6, Qvdow6, Xvdow6, Ewdow6, Lwdow6, Swdow6, Zwdow6;
wire Gxdow6, Nxdow6, Uxdow6, Bydow6, Iydow6, Pydow6, Wydow6, Dzdow6, Kzdow6, Rzdow6;
wire Yzdow6, F0eow6, M0eow6, T0eow6, A1eow6, H1eow6, O1eow6, V1eow6, C2eow6, J2eow6;
wire Q2eow6, X2eow6, E3eow6, L3eow6, S3eow6, Z3eow6, G4eow6, N4eow6, U4eow6, B5eow6;
wire I5eow6, P5eow6, W5eow6, D6eow6, K6eow6, R6eow6, Y6eow6, F7eow6, M7eow6, T7eow6;
wire A8eow6, H8eow6, O8eow6, V8eow6, C9eow6, J9eow6, Q9eow6, X9eow6, Eaeow6, Laeow6;
wire Saeow6, Zaeow6, Gbeow6, Nbeow6, Ubeow6, Bceow6, Iceow6, Pceow6, Wceow6, Ddeow6;
wire Kdeow6, Rdeow6, Ydeow6, Feeow6, Meeow6, Teeow6, Afeow6, Hfeow6, Ofeow6, Vfeow6;
wire Cgeow6, Jgeow6, Qgeow6, Xgeow6, Eheow6, Lheow6, Sheow6, Zheow6, Gieow6, Nieow6;
wire Uieow6, Bjeow6, Ijeow6, Pjeow6, Wjeow6, Dkeow6, Kkeow6, Rkeow6, Ykeow6, Fleow6;
wire Mleow6, Tleow6, Ameow6, Hmeow6, Omeow6, Vmeow6, Cneow6, Jneow6, Qneow6, Xneow6;
wire Eoeow6, Loeow6, Soeow6, Zoeow6, Gpeow6, Npeow6, Upeow6, Bqeow6, Iqeow6, Pqeow6;
wire Wqeow6, Dreow6, Kreow6, Rreow6, Yreow6, Fseow6, Mseow6, Tseow6, Ateow6, Hteow6;
wire Oteow6, Vteow6, Cueow6, Jueow6, Queow6, Xueow6, Eveow6, Lveow6, Sveow6, Zveow6;
wire Gweow6, Nweow6, Uweow6, Bxeow6, Ixeow6, Pxeow6, Wxeow6, Dyeow6, Kyeow6, Ryeow6;
wire Yyeow6, Fzeow6, Mzeow6, Tzeow6, A0fow6, H0fow6, O0fow6, V0fow6, C1fow6, J1fow6;
wire Q1fow6, X1fow6, E2fow6, L2fow6, S2fow6, Z2fow6, G3fow6, N3fow6, U3fow6, B4fow6;
wire I4fow6, P4fow6, W4fow6, D5fow6, K5fow6, R5fow6, Y5fow6, F6fow6, M6fow6, T6fow6;
wire A7fow6, H7fow6, O7fow6, V7fow6, C8fow6, J8fow6, Q8fow6, X8fow6, E9fow6, L9fow6;
wire S9fow6, Z9fow6, Gafow6, Nafow6, Uafow6, Bbfow6, Ibfow6, Pbfow6, Wbfow6, Dcfow6;
wire Kcfow6, Rcfow6, Ycfow6, Fdfow6, Mdfow6, Tdfow6, Aefow6, Hefow6, Oefow6, Vefow6;
wire Cffow6, Jffow6, Qffow6, Xffow6, Egfow6, Lgfow6, Sgfow6, Zgfow6, Ghfow6, Nhfow6;
wire Uhfow6, Bifow6, Iifow6, Pifow6, Wifow6, Djfow6, Kjfow6, Rjfow6, Yjfow6, Fkfow6;
wire Mkfow6, Tkfow6, Alfow6, Hlfow6, Olfow6, Vlfow6, Cmfow6, Jmfow6, Qmfow6, Xmfow6;
wire Enfow6, Lnfow6, Snfow6, Znfow6, Gofow6, Nofow6, Uofow6, Bpfow6, Ipfow6, Ppfow6;
wire Wpfow6, Dqfow6, Kqfow6, Rqfow6, Yqfow6, Frfow6, Mrfow6, Trfow6, Asfow6, Hsfow6;
wire Osfow6, Vsfow6, Ctfow6, Jtfow6, Qtfow6, Xtfow6, Eufow6, Lufow6, Sufow6, Zufow6;
wire Gvfow6, Nvfow6, Uvfow6, Bwfow6, Iwfow6, Pwfow6, Wwfow6, Dxfow6, Kxfow6, Rxfow6;
wire Yxfow6, Fyfow6, Myfow6, Tyfow6, Azfow6, Hzfow6, Ozfow6, Vzfow6, C0gow6, J0gow6;
wire Q0gow6, X0gow6, E1gow6, L1gow6, S1gow6, Z1gow6, G2gow6, N2gow6, U2gow6, B3gow6;
wire I3gow6, P3gow6, W3gow6, D4gow6, K4gow6, R4gow6, Y4gow6, F5gow6, M5gow6, T5gow6;
wire A6gow6, H6gow6, O6gow6, V6gow6, C7gow6, J7gow6, Q7gow6, X7gow6, E8gow6, L8gow6;
wire S8gow6, Z8gow6, G9gow6, N9gow6, U9gow6, Bagow6, Iagow6, Pagow6, Wagow6, Dbgow6;
wire Kbgow6, Rbgow6, Ybgow6, Fcgow6, Mcgow6, Tcgow6, Adgow6, Hdgow6, Odgow6, Vdgow6;
wire Cegow6, Jegow6, Qegow6, Xegow6, Efgow6, Lfgow6, Sfgow6, Zfgow6, Gggow6, Nggow6;
wire Uggow6, Bhgow6, Ihgow6, Phgow6, Whgow6, Digow6, Kigow6, Rigow6, Yigow6, Fjgow6;
wire Mjgow6, Tjgow6, Akgow6, Hkgow6, Okgow6, Vkgow6, Clgow6, Jlgow6, Qlgow6, Xlgow6;
wire Emgow6, Lmgow6, Smgow6, Zmgow6, Gngow6, Nngow6, Ungow6, Bogow6, Iogow6, Pogow6;
wire Wogow6, Dpgow6, Kpgow6, Rpgow6, Ypgow6, Fqgow6, Mqgow6, Tqgow6, Argow6, Hrgow6;
wire Orgow6, Vrgow6, Csgow6, Jsgow6, Qsgow6, Xsgow6, Etgow6, Ltgow6, Stgow6, Ztgow6;
wire Gugow6, Nugow6, Uugow6, Bvgow6, Ivgow6, Pvgow6, Wvgow6, Dwgow6, Kwgow6, Rwgow6;
wire Ywgow6, Fxgow6, Mxgow6, Txgow6, Aygow6, Hygow6, Oygow6, Vygow6, Czgow6, Jzgow6;
wire Qzgow6, Xzgow6, E0how6, L0how6, S0how6, Z0how6, G1how6, N1how6, U1how6, B2how6;
wire I2how6, P2how6, W2how6, D3how6, K3how6, R3how6, Y3how6, F4how6, M4how6, T4how6;
wire A5how6, H5how6, O5how6, V5how6, C6how6, J6how6, Q6how6, X6how6, E7how6, L7how6;
wire S7how6, Z7how6, G8how6, N8how6, U8how6, B9how6, I9how6, P9how6, W9how6, Dahow6;
wire Kahow6, Rahow6, Yahow6, Fbhow6, Mbhow6, Tbhow6, Achow6, Hchow6, Ochow6, Vchow6;
wire Cdhow6, Jdhow6, Qdhow6, Xdhow6, Eehow6, Lehow6, Sehow6, Zehow6, Gfhow6, Nfhow6;
wire Ufhow6, Bghow6, Ighow6, Pghow6, Wghow6, Dhhow6, Khhow6, Rhhow6, Yhhow6, Fihow6;
wire Mihow6, Tihow6, Ajhow6, Hjhow6, Ojhow6, Vjhow6, Ckhow6, Jkhow6, Qkhow6, Xkhow6;
wire Elhow6, Llhow6, Slhow6, Zlhow6, Gmhow6, Nmhow6, Umhow6, Bnhow6, Inhow6, Pnhow6;
wire Wnhow6, Dohow6, Kohow6, Rohow6, Yohow6, Fphow6, Mphow6, Tphow6, Aqhow6, Hqhow6;
wire Oqhow6, Vqhow6, Crhow6, Jrhow6, Qrhow6, Xrhow6, Eshow6, Lshow6, Sshow6, Zshow6;
wire Gthow6, Nthow6, Uthow6, Buhow6, Iuhow6, Puhow6, Wuhow6, Dvhow6, Kvhow6, Rvhow6;
wire Yvhow6, Fwhow6, Mwhow6, Twhow6, Axhow6, Hxhow6, Oxhow6, Vxhow6, Cyhow6, Jyhow6;
wire Qyhow6, Xyhow6, Ezhow6, Lzhow6, Szhow6, Zzhow6, G0iow6, N0iow6, U0iow6, B1iow6;
wire I1iow6, P1iow6, W1iow6, D2iow6, K2iow6, R2iow6, Y2iow6, F3iow6, M3iow6, T3iow6;
wire A4iow6, H4iow6, O4iow6, V4iow6, C5iow6, J5iow6, Q5iow6, X5iow6, E6iow6, L6iow6;
wire S6iow6, Z6iow6, G7iow6, N7iow6, U7iow6, B8iow6, I8iow6, P8iow6, W8iow6, D9iow6;
wire K9iow6, R9iow6, Y9iow6, Faiow6, Maiow6, Taiow6, Abiow6, Hbiow6, Obiow6, Vbiow6;
wire Cciow6, Jciow6, Qciow6, Xciow6, Ediow6, Ldiow6, Sdiow6, Zdiow6, Geiow6, Neiow6;
wire Ueiow6, Bfiow6, Ifiow6, Pfiow6, Wfiow6, Dgiow6, Kgiow6, Rgiow6, Ygiow6, Fhiow6;
wire Mhiow6, Thiow6, Aiiow6, Hiiow6, Oiiow6, Viiow6, Cjiow6, Jjiow6, Qjiow6, Xjiow6;
wire Ekiow6, Lkiow6, Skiow6, Zkiow6, Gliow6, Nliow6, Uliow6, Bmiow6, Imiow6, Pmiow6;
wire Wmiow6, Dniow6, Kniow6, Rniow6, Yniow6, Foiow6, Moiow6, Toiow6, Apiow6, Hpiow6;
wire Opiow6, Vpiow6, Cqiow6, Jqiow6, Qqiow6, Xqiow6, Eriow6, Lriow6, Sriow6, Zriow6;
wire Gsiow6, Nsiow6, Usiow6, Btiow6, Itiow6, Ptiow6, Wtiow6, Duiow6, Kuiow6, Ruiow6;
wire Yuiow6, Fviow6, Mviow6, Tviow6, Awiow6, Hwiow6, Owiow6, Vwiow6, Cxiow6, Jxiow6;
wire Qxiow6, Xxiow6, Eyiow6, Lyiow6, Syiow6, Zyiow6, Gziow6, Nziow6, Uziow6, B0jow6;
wire I0jow6, P0jow6, W0jow6, D1jow6, K1jow6, R1jow6, Y1jow6, F2jow6, M2jow6, T2jow6;
wire A3jow6, H3jow6, O3jow6, V3jow6, C4jow6, J4jow6, Q4jow6, X4jow6, E5jow6, L5jow6;
wire S5jow6, Z5jow6, G6jow6, N6jow6, U6jow6, B7jow6, I7jow6, P7jow6, W7jow6, D8jow6;
wire K8jow6, R8jow6, Y8jow6, F9jow6, M9jow6, T9jow6, Aajow6, Hajow6, Oajow6, Vajow6;
wire Cbjow6, Jbjow6, Qbjow6, Xbjow6, Ecjow6, Lcjow6, Scjow6, Zcjow6, Gdjow6, Ndjow6;
wire Udjow6, Bejow6, Iejow6, Pejow6, Wejow6, Dfjow6, Kfjow6, Rfjow6, Yfjow6, Fgjow6;
wire Mgjow6, Tgjow6, Ahjow6, Hhjow6, Ohjow6, Vhjow6, Cijow6, Jijow6, Qijow6, Xijow6;
wire Ejjow6, Ljjow6, Sjjow6, Zjjow6, Gkjow6, Nkjow6, Ukjow6, Bljow6, Iljow6, Pljow6;
wire Wljow6, Dmjow6, Kmjow6, Rmjow6, Ymjow6, Fnjow6, Mnjow6, Tnjow6, Aojow6, Hojow6;
wire Oojow6, Vojow6, Cpjow6, Jpjow6, Qpjow6, Xpjow6, Eqjow6, Lqjow6, Sqjow6, Zqjow6;
wire Grjow6, Nrjow6, Urjow6, Bsjow6, Isjow6, Psjow6, Wsjow6, Dtjow6, Ktjow6, Rtjow6;
wire Ytjow6, Fujow6, Mujow6, Tujow6, Avjow6, Hvjow6, Ovjow6, Vvjow6, Cwjow6, Jwjow6;
wire Qwjow6, Xwjow6, Exjow6, Lxjow6, Sxjow6, Zxjow6, Gyjow6, Nyjow6, Uyjow6, Bzjow6;
wire Izjow6, Pzjow6, Wzjow6, D0kow6, K0kow6, R0kow6, Y0kow6, F1kow6, M1kow6, T1kow6;
wire A2kow6, H2kow6, O2kow6, V2kow6, C3kow6, J3kow6, Q3kow6, X3kow6, E4kow6, L4kow6;
wire S4kow6, Z4kow6, G5kow6, N5kow6, U5kow6, B6kow6, I6kow6, P6kow6, W6kow6, D7kow6;
wire K7kow6, R7kow6, Y7kow6, F8kow6, M8kow6, T8kow6, A9kow6, H9kow6, O9kow6, V9kow6;
wire Cakow6, Jakow6, Qakow6, Xakow6, Ebkow6, Lbkow6, Sbkow6, Zbkow6, Gckow6, Nckow6;
wire Uckow6, Bdkow6, Idkow6, Pdkow6, Wdkow6, Dekow6, Kekow6, Rekow6, Yekow6, Ffkow6;
wire Mfkow6, Tfkow6, Agkow6, Hgkow6, Ogkow6, Vgkow6, Chkow6, Jhkow6, Qhkow6, Xhkow6;
wire Eikow6, Likow6, Sikow6, Zikow6, Gjkow6, Njkow6, Ujkow6, Bkkow6, Ikkow6, Pkkow6;
wire Wkkow6, Dlkow6, Klkow6, Rlkow6, Ylkow6, Fmkow6, Mmkow6, Tmkow6, Ankow6, Hnkow6;
wire Onkow6, Vnkow6, Cokow6, Jokow6, Qokow6, Xokow6, Epkow6, Lpkow6, Spkow6, Zpkow6;
wire Gqkow6, Nqkow6, Uqkow6, Brkow6, Irkow6, Prkow6, Wrkow6, Dskow6, Kskow6, Rskow6;
wire Yskow6, Ftkow6, Mtkow6, Ttkow6, Aukow6, Hukow6, Oukow6, Vukow6, Cvkow6, Jvkow6;
wire Qvkow6, Xvkow6, Ewkow6, Lwkow6, Swkow6, Zwkow6, Gxkow6, Nxkow6, Uxkow6, Bykow6;
wire Iykow6, Pykow6, Wykow6, Dzkow6, Kzkow6, Rzkow6, Yzkow6, F0low6, M0low6, T0low6;
wire A1low6, H1low6, O1low6, V1low6, C2low6, J2low6, Q2low6, X2low6, E3low6, L3low6;
wire S3low6, Z3low6, G4low6, N4low6, U4low6, B5low6, I5low6, P5low6, W5low6, D6low6;
wire K6low6, R6low6, Y6low6, F7low6, M7low6, T7low6, A8low6, H8low6, O8low6, V8low6;
wire C9low6, J9low6, Q9low6, X9low6, Ealow6, Lalow6, Salow6, Zalow6, Gblow6, Nblow6;
wire Ublow6, Bclow6, Iclow6, Pclow6, Wclow6, Ddlow6, Kdlow6, Rdlow6, Ydlow6, Felow6;
wire Melow6, Telow6, Aflow6, Hflow6, Oflow6, Vflow6, Cglow6, Jglow6, Qglow6, Xglow6;
wire Ehlow6, Lhlow6, Shlow6, Zhlow6, Gilow6, Nilow6, Uilow6, Bjlow6, Ijlow6, Pjlow6;
wire Wjlow6, Dklow6, Kklow6, Rklow6, Yklow6, Fllow6, Mllow6, Tllow6, Amlow6, Hmlow6;
wire Omlow6, Vmlow6, Cnlow6, Jnlow6, Qnlow6, Xnlow6, Eolow6, Lolow6, Solow6, Zolow6;
wire Gplow6, Nplow6, Uplow6, Bqlow6, Iqlow6, Pqlow6, Wqlow6, Drlow6, Krlow6, Rrlow6;
wire Yrlow6, Fslow6, Mslow6, Tslow6, Atlow6, Htlow6, Otlow6, Vtlow6, Culow6, Julow6;
wire Qulow6, Xulow6, Evlow6, Lvlow6, Svlow6, Zvlow6, Gwlow6, Nwlow6, Uwlow6, Bxlow6;
wire Ixlow6, Pxlow6, Wxlow6, Dylow6, Kylow6, Rylow6, Yylow6, Fzlow6, Mzlow6, Tzlow6;
wire A0mow6, H0mow6, O0mow6, V0mow6, C1mow6, J1mow6, Q1mow6, X1mow6, E2mow6, L2mow6;
wire S2mow6, Z2mow6, G3mow6, N3mow6, U3mow6, B4mow6, I4mow6, P4mow6, W4mow6, D5mow6;
wire K5mow6, R5mow6, Y5mow6, F6mow6, M6mow6, T6mow6, A7mow6, H7mow6, O7mow6, V7mow6;
wire C8mow6, J8mow6, Q8mow6, X8mow6, E9mow6, L9mow6, S9mow6, Z9mow6, Gamow6, Namow6;
wire Uamow6, Bbmow6, Ibmow6, Pbmow6, Wbmow6, Dcmow6, Kcmow6, Rcmow6, Ycmow6, Fdmow6;
wire Mdmow6, Tdmow6, Aemow6, Hemow6, Oemow6, Vemow6, Cfmow6, Jfmow6, Qfmow6, Xfmow6;
wire Egmow6, Lgmow6, Sgmow6, Zgmow6, Ghmow6, Nhmow6, Uhmow6, Bimow6, Iimow6, Pimow6;
wire Wimow6, Djmow6, Kjmow6, Rjmow6, Yjmow6, Fkmow6, Mkmow6, Tkmow6, Almow6, Hlmow6;
wire Olmow6, Vlmow6, Cmmow6, Jmmow6, Qmmow6, Xmmow6, Enmow6, Lnmow6, Snmow6, Znmow6;
wire Gomow6, Nomow6, Uomow6, Bpmow6, Ipmow6, Ppmow6, Wpmow6, Dqmow6, Kqmow6, Rqmow6;
wire Yqmow6, Frmow6, Mrmow6, Trmow6, Asmow6, Hsmow6, Osmow6, Vsmow6, Ctmow6, Jtmow6;
wire Qtmow6, Xtmow6, Eumow6, Lumow6, Sumow6, Zumow6, Gvmow6, Nvmow6, Uvmow6, Bwmow6;
wire Iwmow6, Pwmow6, Wwmow6, Dxmow6, Kxmow6, Rxmow6, Yxmow6, Fymow6, Mymow6, Tymow6;
wire Azmow6, Hzmow6, Ozmow6, Vzmow6, C0now6, J0now6, Q0now6, X0now6, E1now6, L1now6;
wire S1now6, Z1now6, G2now6, N2now6, U2now6, B3now6, I3now6, P3now6, W3now6, D4now6;
wire K4now6, R4now6, Y4now6, F5now6, M5now6, T5now6, A6now6, H6now6, O6now6, V6now6;
wire C7now6, J7now6, Q7now6, X7now6, E8now6, L8now6, S8now6, Z8now6, G9now6, N9now6;
wire U9now6, Banow6, Ianow6, Panow6, Wanow6, Dbnow6, Kbnow6, Rbnow6, Ybnow6, Fcnow6;
wire Mcnow6, Tcnow6, Adnow6, Hdnow6, Odnow6, Vdnow6, Cenow6, Jenow6, Qenow6, Xenow6;
wire Efnow6, Lfnow6, Sfnow6, Zfnow6, Ggnow6, Ngnow6, Ugnow6, Bhnow6, Ihnow6, Phnow6;
wire Whnow6, Dinow6, Kinow6, Rinow6, Yinow6, Fjnow6, Mjnow6, Tjnow6, Aknow6, Hknow6;
wire Oknow6, Vknow6, Clnow6, Jlnow6, Qlnow6, Xlnow6, Emnow6, Lmnow6, Smnow6, Zmnow6;
wire Gnnow6, Nnnow6, Unnow6, Bonow6, Ionow6, Ponow6, Wonow6, Dpnow6, Kpnow6, Rpnow6;
wire Ypnow6, Fqnow6, Mqnow6, Tqnow6, Arnow6, Hrnow6, Ornow6, Vrnow6, Csnow6, Jsnow6;
wire Qsnow6, Xsnow6, Etnow6, Ltnow6, Stnow6, Ztnow6, Gunow6, Nunow6, Uunow6, Bvnow6;
wire Ivnow6, Pvnow6, Wvnow6, Dwnow6, Kwnow6, Rwnow6, Ywnow6, Fxnow6, Mxnow6, Txnow6;
wire Aynow6, Hynow6, Oynow6, Vynow6, Cznow6, Jznow6, Qznow6, Xznow6, E0oow6, L0oow6;
wire S0oow6, Z0oow6, G1oow6, N1oow6, U1oow6, B2oow6, I2oow6, P2oow6, W2oow6, D3oow6;
wire K3oow6, R3oow6, Y3oow6, F4oow6, M4oow6, T4oow6, A5oow6, H5oow6, O5oow6, V5oow6;
wire C6oow6, J6oow6, Q6oow6, X6oow6, E7oow6, L7oow6, S7oow6, Z7oow6, G8oow6, N8oow6;
wire U8oow6, B9oow6, I9oow6, P9oow6, W9oow6, Daoow6, Kaoow6, Raoow6, Yaoow6, Fboow6;
wire Mboow6, Tboow6, Acoow6, Hcoow6, Ocoow6, Vcoow6, Cdoow6, Jdoow6, Qdoow6, Xdoow6;
wire Eeoow6, Leoow6, Seoow6, Zeoow6, Gfoow6, Nfoow6, Ufoow6, Bgoow6, Igoow6, Pgoow6;
wire Wgoow6, Dhoow6, Khoow6, Rhoow6, Yhoow6, Fioow6, Mioow6, Tioow6, Ajoow6, Hjoow6;
wire Ojoow6, Vjoow6, Ckoow6, Jkoow6, Qkoow6, Xkoow6, Eloow6, Lloow6, Sloow6, Zloow6;
wire Gmoow6, Nmoow6, Umoow6, Bnoow6, Inoow6, Pnoow6, Wnoow6, Dooow6, Kooow6, Rooow6;
wire Yooow6, Fpoow6, Mpoow6, Tpoow6, Aqoow6, Hqoow6, Oqoow6, Vqoow6, Croow6, Jroow6;
wire Qroow6, Xroow6, Esoow6, Lsoow6, Ssoow6, Zsoow6, Gtoow6, Ntoow6, Utoow6, Buoow6;
wire Iuoow6, Puoow6, Wuoow6, Dvoow6, Kvoow6, Rvoow6, Yvoow6, Fwoow6, Mwoow6, Twoow6;
wire Axoow6, Hxoow6, Oxoow6, Vxoow6, Cyoow6, Jyoow6, Qyoow6, Xyoow6, Ezoow6, Lzoow6;
wire Szoow6, Zzoow6, G0pow6, N0pow6, U0pow6, B1pow6, I1pow6, P1pow6, W1pow6, D2pow6;
wire K2pow6, R2pow6, Y2pow6, F3pow6, M3pow6, T3pow6, A4pow6, H4pow6, O4pow6, V4pow6;
wire C5pow6, J5pow6, Q5pow6, X5pow6, E6pow6, L6pow6, S6pow6, Z6pow6, G7pow6, N7pow6;
wire U7pow6, B8pow6, I8pow6, P8pow6, W8pow6, D9pow6, K9pow6, R9pow6, Y9pow6, Fapow6;
wire Mapow6, Tapow6, Abpow6, Hbpow6, Obpow6, Vbpow6, Ccpow6, Jcpow6, Qcpow6, Xcpow6;
wire Edpow6, Ldpow6, Sdpow6, Zdpow6, Gepow6, Nepow6, Uepow6, Bfpow6, Ifpow6, Pfpow6;
wire Wfpow6, Dgpow6, Kgpow6, Rgpow6, Ygpow6, Fhpow6, Mhpow6, Thpow6, Aipow6, Hipow6;
wire Oipow6, Vipow6, Cjpow6, Jjpow6, Qjpow6, Xjpow6, Ekpow6, Lkpow6, Skpow6, Zkpow6;
wire Glpow6, Nlpow6, Ulpow6, Bmpow6, Impow6, Pmpow6, Wmpow6, Dnpow6, Knpow6, Rnpow6;
wire Ynpow6, Fopow6, Mopow6, Topow6, Appow6, Hppow6, Oppow6, Vppow6, Cqpow6, Jqpow6;
wire Qqpow6, Xqpow6, Erpow6, Lrpow6, Srpow6, Zrpow6, Gspow6, Nspow6, Uspow6, Btpow6;
wire Itpow6, Ptpow6, Wtpow6, Dupow6, Kupow6, Rupow6, Yupow6, Fvpow6, Mvpow6, Tvpow6;
wire Awpow6, Hwpow6, Owpow6, Vwpow6, Cxpow6, Jxpow6, Qxpow6, Xxpow6, Eypow6, Lypow6;
wire Sypow6, Zypow6, Gzpow6, Nzpow6, Uzpow6, B0qow6, I0qow6, P0qow6, W0qow6, D1qow6;
wire K1qow6, R1qow6, Y1qow6, F2qow6, M2qow6, T2qow6, A3qow6, H3qow6, O3qow6, V3qow6;
wire C4qow6, J4qow6, Q4qow6, X4qow6, E5qow6, L5qow6, S5qow6, Z5qow6, G6qow6, N6qow6;
wire U6qow6, B7qow6, I7qow6, P7qow6, W7qow6, D8qow6, K8qow6, R8qow6, Y8qow6, F9qow6;
wire M9qow6, T9qow6, Aaqow6, Haqow6, Oaqow6, Vaqow6, Cbqow6, Jbqow6, Qbqow6, Xbqow6;
wire Ecqow6, Lcqow6, Scqow6, Zcqow6, Gdqow6, Ndqow6, Udqow6, Beqow6, Ieqow6, Peqow6;
wire Weqow6, Dfqow6, Kfqow6, Rfqow6, Yfqow6, Fgqow6, Mgqow6, Tgqow6, Ahqow6, Hhqow6;
wire Ohqow6, Vhqow6, Ciqow6, Jiqow6, Qiqow6, Xiqow6, Ejqow6, Ljqow6, Sjqow6, Zjqow6;
wire Gkqow6, Nkqow6, Ukqow6, Blqow6, Ilqow6, Plqow6, Wlqow6, Dmqow6, Kmqow6, Rmqow6;
wire Ymqow6, Fnqow6, Mnqow6, Tnqow6, Aoqow6, Hoqow6, Ooqow6, Voqow6, Cpqow6, Jpqow6;
wire Qpqow6, Xpqow6, Eqqow6, Lqqow6, Sqqow6, Zqqow6, Grqow6, Nrqow6, Urqow6, Bsqow6;
wire Isqow6, Psqow6, Wsqow6, Dtqow6, Ktqow6, Rtqow6, Ytqow6, Fuqow6, Muqow6, Tuqow6;
wire Avqow6, Hvqow6, Ovqow6, Vvqow6, Cwqow6, Jwqow6, Qwqow6, Xwqow6, Exqow6, Lxqow6;
wire Sxqow6, Zxqow6, Gyqow6, Nyqow6, Uyqow6, Bzqow6, Izqow6, Pzqow6, Wzqow6, D0row6;
wire K0row6, R0row6, Y0row6, F1row6, M1row6, T1row6, A2row6, H2row6, O2row6, V2row6;
wire C3row6, J3row6, Q3row6, X3row6, E4row6, L4row6, S4row6, Z4row6, G5row6, N5row6;
wire U5row6, B6row6, I6row6, P6row6, W6row6, D7row6, K7row6, R7row6, Y7row6, F8row6;
wire M8row6, T8row6, A9row6, H9row6, O9row6, V9row6, Carow6, Jarow6, Qarow6, Xarow6;
wire Ebrow6, Lbrow6, Sbrow6, Zbrow6, Gcrow6, Ncrow6, Ucrow6, Bdrow6, Idrow6, Pdrow6;
wire Wdrow6, Derow6, Kerow6, Rerow6, Yerow6, Ffrow6, Mfrow6, Tfrow6, Agrow6, Hgrow6;
wire Ogrow6, Vgrow6, Chrow6, Jhrow6, Qhrow6, Xhrow6, Eirow6, Lirow6, Sirow6, Zirow6;
wire Gjrow6, Njrow6, Ujrow6, Bkrow6, Ikrow6, Pkrow6, Wkrow6, Dlrow6, Klrow6, Rlrow6;
wire Ylrow6, Fmrow6, Mmrow6, Tmrow6, Anrow6, Hnrow6, Onrow6, Vnrow6, Corow6, Jorow6;
wire Qorow6, Xorow6, Eprow6, Lprow6, Sprow6, Zprow6, Gqrow6, Nqrow6, Uqrow6, Brrow6;
wire Irrow6, Prrow6, Wrrow6, Dsrow6, Ksrow6, Rsrow6, Ysrow6, Ftrow6, Mtrow6, Ttrow6;
wire Aurow6, Hurow6, Ourow6, Vurow6, Cvrow6, Jvrow6, Qvrow6, Xvrow6, Ewrow6, Lwrow6;
wire Swrow6, Zwrow6, Gxrow6, Nxrow6, Uxrow6, Byrow6, Iyrow6, Pyrow6, Wyrow6, Dzrow6;
wire Kzrow6, Rzrow6, Yzrow6, F0sow6, M0sow6, T0sow6, A1sow6, H1sow6, O1sow6, V1sow6;
wire C2sow6, J2sow6, Q2sow6, X2sow6, E3sow6, L3sow6, S3sow6, Z3sow6, G4sow6, N4sow6;
wire U4sow6, B5sow6, I5sow6, P5sow6, W5sow6, D6sow6, K6sow6, R6sow6, Y6sow6, F7sow6;
wire M7sow6, T7sow6, A8sow6, H8sow6, O8sow6, V8sow6, C9sow6, J9sow6, Q9sow6, X9sow6;
wire Easow6, Lasow6, Sasow6, Zasow6, Gbsow6, Nbsow6, Ubsow6, Bcsow6, Icsow6, Pcsow6;
wire Wcsow6, Ddsow6, Kdsow6, Rdsow6, Ydsow6, Fesow6, Mesow6, Tesow6, Afsow6, Hfsow6;
wire Ofsow6, Vfsow6, Cgsow6, Jgsow6, Qgsow6, Xgsow6, Ehsow6, Lhsow6, Shsow6, Zhsow6;
wire Gisow6, Nisow6, Uisow6, Bjsow6, Ijsow6, Pjsow6, Wjsow6, Dksow6, Kksow6, Rksow6;
wire Yksow6, Flsow6, Mlsow6, Tlsow6, Amsow6, Hmsow6, Omsow6, Vmsow6, Cnsow6, Jnsow6;
wire Qnsow6, Xnsow6, Eosow6, Losow6, Sosow6, Zosow6, Gpsow6, Npsow6, Upsow6, Bqsow6;
wire Iqsow6, Pqsow6, Wqsow6, Drsow6, Krsow6, Rrsow6, Yrsow6, Fssow6, Mssow6, Tssow6;
wire Atsow6, Htsow6, Otsow6, Vtsow6, Cusow6, Jusow6, Qusow6, Xusow6, Evsow6, Lvsow6;
wire Svsow6, Zvsow6, Gwsow6, Nwsow6, Uwsow6, Bxsow6, Ixsow6, Pxsow6, Wxsow6, Dysow6;
wire Kysow6, Rysow6, Yysow6, Fzsow6, Mzsow6, Tzsow6, A0tow6, H0tow6, O0tow6, V0tow6;
wire C1tow6, J1tow6, Q1tow6, X1tow6, E2tow6, L2tow6, S2tow6, Z2tow6, G3tow6, N3tow6;
wire U3tow6, B4tow6, I4tow6, P4tow6, W4tow6, D5tow6, K5tow6, R5tow6, Y5tow6, F6tow6;
wire M6tow6, T6tow6, A7tow6, H7tow6, O7tow6, V7tow6, C8tow6, J8tow6, Q8tow6, X8tow6;
wire E9tow6, L9tow6, S9tow6, Z9tow6, Gatow6, Natow6, Uatow6, Bbtow6, Ibtow6, Pbtow6;
wire Wbtow6, Dctow6, Kctow6, Rctow6, Yctow6, Fdtow6, Mdtow6, Tdtow6, Aetow6, Hetow6;
wire Oetow6, Vetow6, Cftow6, Jftow6, Qftow6, Xftow6, Egtow6, Lgtow6, Sgtow6, Zgtow6;
wire Ghtow6, Nhtow6, Uhtow6, Bitow6, Iitow6, Pitow6, Witow6, Djtow6, Kjtow6, Rjtow6;
wire Yjtow6, Fktow6, Mktow6, Tktow6, Altow6, Hltow6, Oltow6, Vltow6, Cmtow6, Jmtow6;
wire Qmtow6, Xmtow6, Entow6, Lntow6, Sntow6, Zntow6, Gotow6, Notow6, Uotow6, Bptow6;
wire Iptow6, Pptow6, Wptow6, Dqtow6, Kqtow6, Rqtow6, Yqtow6, Frtow6, Mrtow6, Trtow6;
wire Astow6, Hstow6, Ostow6, Vstow6, Cttow6, Jttow6, Qttow6, Xttow6, Eutow6, Lutow6;
wire Sutow6, Zutow6, Gvtow6, Nvtow6, Uvtow6, Bwtow6, Iwtow6, Pwtow6, Wwtow6, Dxtow6;
wire Kxtow6, Rxtow6, Yxtow6, Fytow6, Mytow6, Tytow6, Aztow6, Hztow6, Oztow6, Vztow6;
wire C0uow6, J0uow6, Q0uow6, X0uow6, E1uow6, L1uow6, S1uow6, Z1uow6, G2uow6, N2uow6;
wire U2uow6, B3uow6, I3uow6, P3uow6, W3uow6, D4uow6, K4uow6, R4uow6, Y4uow6, F5uow6;
wire M5uow6, T5uow6, A6uow6, H6uow6, O6uow6, V6uow6, C7uow6, J7uow6, Q7uow6, X7uow6;
wire E8uow6, L8uow6, S8uow6, Z8uow6, G9uow6, N9uow6, U9uow6, Bauow6, Iauow6, Pauow6;
wire Wauow6, Dbuow6, Kbuow6, Rbuow6, Ybuow6, Fcuow6, Mcuow6, Tcuow6, Aduow6, Hduow6;
wire Oduow6, Vduow6, Ceuow6, Jeuow6, Qeuow6, Xeuow6, Efuow6, Lfuow6, Sfuow6, Zfuow6;
wire Gguow6, Nguow6, Uguow6, Bhuow6, Ihuow6, Phuow6, Whuow6, Diuow6, Kiuow6, Riuow6;
wire Yiuow6, Fjuow6, Mjuow6, Tjuow6, Akuow6, Hkuow6, Okuow6, Vkuow6, Cluow6, Jluow6;
wire Qluow6, Xluow6, Emuow6, Lmuow6, Smuow6, Zmuow6, Gnuow6, Nnuow6, Unuow6, Bouow6;
wire Iouow6, Pouow6, Wouow6, Dpuow6, Kpuow6, Rpuow6, Ypuow6, Fquow6, Mquow6, Tquow6;
wire Aruow6, Hruow6, Oruow6, Vruow6, Csuow6, Jsuow6, Qsuow6, Xsuow6, Etuow6, Ltuow6;
wire Stuow6, Ztuow6, Guuow6, Nuuow6, Uuuow6, Bvuow6, Ivuow6, Pvuow6, Wvuow6, Dwuow6;
wire Kwuow6, Rwuow6, Ywuow6, Fxuow6, Mxuow6, Txuow6, Ayuow6, Hyuow6, Oyuow6, Vyuow6;
wire Czuow6, Jzuow6, Qzuow6, Xzuow6, E0vow6, L0vow6, S0vow6, Z0vow6, G1vow6, N1vow6;
wire U1vow6, B2vow6, I2vow6, P2vow6, W2vow6, D3vow6, K3vow6, R3vow6, Y3vow6, F4vow6;
wire M4vow6, T4vow6, A5vow6, H5vow6, O5vow6, V5vow6, C6vow6, J6vow6, Q6vow6, X6vow6;
wire E7vow6, L7vow6, S7vow6, Z7vow6, G8vow6, N8vow6, U8vow6, B9vow6, I9vow6, P9vow6;
wire W9vow6, Davow6, Kavow6, Ravow6, Yavow6, Fbvow6, Mbvow6, Tbvow6, Acvow6, Hcvow6;
wire Ocvow6, Vcvow6, Cdvow6, Jdvow6, Qdvow6, Xdvow6, Eevow6, Levow6, Sevow6, Zevow6;
wire Gfvow6, Nfvow6, Ufvow6, Bgvow6, Igvow6, Pgvow6, Wgvow6, Dhvow6, Khvow6, Rhvow6;
wire Yhvow6, Fivow6, Mivow6, Tivow6, Ajvow6, Hjvow6, Ojvow6, Vjvow6, Ckvow6, Jkvow6;
wire Qkvow6, Xkvow6, Elvow6, Llvow6, Slvow6, Zlvow6, Gmvow6, Nmvow6, Umvow6, Bnvow6;
wire Invow6, Pnvow6, Wnvow6, Dovow6, Kovow6, Rovow6, Yovow6, Fpvow6, Mpvow6, Tpvow6;
wire Aqvow6, Hqvow6, Oqvow6, Vqvow6, Crvow6, Jrvow6, Qrvow6, Xrvow6, Esvow6, Lsvow6;
wire Ssvow6, Zsvow6, Gtvow6, Ntvow6, Utvow6, Buvow6, Iuvow6, Puvow6, Wuvow6, Dvvow6;
wire Kvvow6, Rvvow6, Yvvow6, Fwvow6, Mwvow6, Twvow6, Axvow6, Hxvow6, Oxvow6, Vxvow6;
wire Cyvow6, Jyvow6, Qyvow6, Xyvow6, Ezvow6, Lzvow6, Szvow6, Zzvow6, G0wow6, N0wow6;
wire U0wow6, B1wow6, I1wow6, P1wow6, W1wow6, D2wow6, K2wow6, R2wow6, Y2wow6, F3wow6;
wire M3wow6, T3wow6, A4wow6, H4wow6, O4wow6, V4wow6, C5wow6, J5wow6, Q5wow6, X5wow6;
wire E6wow6, L6wow6, S6wow6, Z6wow6, G7wow6, N7wow6, U7wow6, B8wow6, I8wow6, P8wow6;
wire W8wow6, D9wow6, K9wow6, R9wow6, Y9wow6, Fawow6, Mawow6, Tawow6, Abwow6, Hbwow6;
wire Obwow6, Vbwow6, Ccwow6, Jcwow6, Qcwow6, Xcwow6, Edwow6, Ldwow6, Sdwow6, Zdwow6;
wire Gewow6, Newow6, Uewow6, Bfwow6, Ifwow6, Pfwow6, Wfwow6, Dgwow6, Kgwow6, Rgwow6;
wire Ygwow6, Fhwow6, Mhwow6, Thwow6, Aiwow6, Hiwow6, Oiwow6, Viwow6, Cjwow6, Jjwow6;
wire Qjwow6, Xjwow6, Ekwow6, Lkwow6, Skwow6, Zkwow6, Glwow6, Nlwow6, Ulwow6, Bmwow6;
wire Imwow6, Pmwow6, Wmwow6, Dnwow6, Knwow6, Rnwow6, Ynwow6, Fowow6, Mowow6, Towow6;
wire Apwow6, Hpwow6, Opwow6, Vpwow6, Cqwow6, Jqwow6, Qqwow6, Xqwow6, Erwow6, Lrwow6;
wire Srwow6, Zrwow6, Gswow6, Nswow6, Uswow6, Btwow6, Itwow6, Ptwow6, Wtwow6, Duwow6;
wire Kuwow6, Ruwow6, Yuwow6, Fvwow6, Mvwow6, Tvwow6, Awwow6, Hwwow6, Owwow6, Vwwow6;
wire Cxwow6, Jxwow6, Qxwow6, Xxwow6, Eywow6, Lywow6, Sywow6, Zywow6, Gzwow6, Nzwow6;
wire Uzwow6, B0xow6, I0xow6, P0xow6, W0xow6, D1xow6, K1xow6, R1xow6, Y1xow6, F2xow6;
wire M2xow6, T2xow6, A3xow6, H3xow6, O3xow6, V3xow6, C4xow6, J4xow6, Q4xow6, X4xow6;
wire E5xow6, L5xow6, S5xow6, Z5xow6, G6xow6, N6xow6, U6xow6, B7xow6, I7xow6, P7xow6;
wire W7xow6, D8xow6, K8xow6, R8xow6, Y8xow6, F9xow6, M9xow6, T9xow6, Aaxow6, Haxow6;
wire Oaxow6, Vaxow6, Cbxow6, Jbxow6, Qbxow6, Xbxow6, Ecxow6, Lcxow6, Scxow6, Zcxow6;
wire Gdxow6, Ndxow6, Udxow6, Bexow6, Iexow6, Pexow6, Wexow6, Dfxow6, Kfxow6, Rfxow6;
wire Yfxow6, Fgxow6, Mgxow6, Tgxow6, Ahxow6, Hhxow6, Ohxow6, Vhxow6, Cixow6, Jixow6;
wire Qixow6, Xixow6, Ejxow6, Ljxow6, Sjxow6, Zjxow6, Gkxow6, Nkxow6, Ukxow6, Blxow6;
wire Ilxow6, Plxow6, Wlxow6, Dmxow6, Kmxow6, Rmxow6, Ymxow6, Fnxow6, Mnxow6, Tnxow6;
wire Aoxow6, Hoxow6, Ooxow6, Voxow6, Cpxow6, Jpxow6, Qpxow6, Xpxow6, Eqxow6, Lqxow6;
wire Sqxow6, Zqxow6, Grxow6, Nrxow6, Urxow6, Bsxow6, Isxow6, Psxow6, Wsxow6, Dtxow6;
wire Ktxow6, Rtxow6, Ytxow6, Fuxow6, Muxow6, Tuxow6, Avxow6, Hvxow6, Ovxow6, Vvxow6;
wire Cwxow6, Jwxow6, Qwxow6, Xwxow6, Exxow6, Lxxow6, Sxxow6, Zxxow6, Gyxow6, Nyxow6;
wire Uyxow6, Bzxow6, Izxow6, Pzxow6, Wzxow6, D0yow6, K0yow6, R0yow6, Y0yow6, F1yow6;
wire M1yow6, T1yow6, A2yow6, H2yow6, O2yow6, V2yow6, C3yow6, J3yow6, Q3yow6, X3yow6;
wire E4yow6, L4yow6, S4yow6, Z4yow6, G5yow6, N5yow6, U5yow6, B6yow6, I6yow6, P6yow6;
wire W6yow6, D7yow6, K7yow6, R7yow6, Y7yow6, F8yow6, M8yow6, T8yow6, A9yow6, H9yow6;
wire O9yow6, V9yow6, Cayow6, Jayow6, Qayow6, Xayow6, Ebyow6, Lbyow6, Sbyow6, Zbyow6;
wire Gcyow6, Ncyow6, Ucyow6, Bdyow6, Idyow6, Pdyow6, Wdyow6, Deyow6, Keyow6, Reyow6;
wire Yeyow6, Ffyow6, Mfyow6, Tfyow6, Agyow6, Hgyow6, Ogyow6, Vgyow6, Chyow6, Jhyow6;
wire Qhyow6, Xhyow6, Eiyow6, Liyow6, Siyow6, Ziyow6, Gjyow6, Njyow6, Ujyow6, Bkyow6;
wire Ikyow6, Pkyow6, Wkyow6, Dlyow6, Klyow6, Rlyow6, Ylyow6, Fmyow6, Mmyow6, Tmyow6;
wire Anyow6, Hnyow6, Onyow6, Vnyow6, Coyow6, Joyow6, Qoyow6, Xoyow6, Epyow6, Lpyow6;
wire Spyow6, Zpyow6, Gqyow6, Nqyow6, Uqyow6, Bryow6, Iryow6, Pryow6, Wryow6, Dsyow6;
wire Ksyow6, Rsyow6, Ysyow6, Ftyow6, Mtyow6, Ttyow6, Auyow6, Huyow6, Ouyow6, Vuyow6;
wire Cvyow6, Jvyow6, Qvyow6, Xvyow6, Ewyow6, Lwyow6, Swyow6, Zwyow6, Gxyow6, Nxyow6;
wire Uxyow6, Byyow6, Iyyow6, Pyyow6, Wyyow6, Dzyow6, Kzyow6, Rzyow6, Yzyow6, F0zow6;
wire M0zow6, T0zow6, A1zow6, H1zow6, O1zow6, V1zow6, C2zow6, J2zow6, Q2zow6, X2zow6;
wire E3zow6, L3zow6, S3zow6, Z3zow6, G4zow6, N4zow6, U4zow6, B5zow6, I5zow6, P5zow6;
wire W5zow6, D6zow6, K6zow6, R6zow6, Y6zow6, F7zow6, M7zow6, T7zow6, A8zow6, H8zow6;
wire O8zow6, V8zow6, C9zow6, J9zow6, Q9zow6, X9zow6, Eazow6, Lazow6, Sazow6, Zazow6;
wire Gbzow6, Nbzow6, Ubzow6, Bczow6, Iczow6, Pczow6, Wczow6, Ddzow6, Kdzow6, Rdzow6;
wire Ydzow6, Fezow6, Mezow6, Tezow6, Afzow6, Hfzow6, Ofzow6, Vfzow6, Cgzow6, Jgzow6;
wire Qgzow6, Xgzow6, Ehzow6, Lhzow6, Shzow6, Zhzow6, Gizow6, Nizow6, Uizow6, Bjzow6;
wire Ijzow6, Pjzow6, Wjzow6, Dkzow6, Kkzow6, Rkzow6, Ykzow6, Flzow6, Mlzow6, Tlzow6;
wire Amzow6, Hmzow6, Omzow6, Vmzow6, Cnzow6, Jnzow6, Qnzow6, Xnzow6, Eozow6, Lozow6;
wire Sozow6, Zozow6, Gpzow6, Npzow6, Upzow6, Bqzow6, Iqzow6, Pqzow6, Wqzow6, Drzow6;
wire Krzow6, Rrzow6, Yrzow6, Fszow6, Mszow6, Tszow6, Atzow6, Htzow6, Otzow6, Vtzow6;
wire Cuzow6, Juzow6, Quzow6, Xuzow6, Evzow6, Lvzow6, Svzow6, Zvzow6, Gwzow6, Nwzow6;
wire Uwzow6, Bxzow6, Ixzow6, Pxzow6, Wxzow6, Dyzow6, Kyzow6, Ryzow6, Yyzow6, Fzzow6;
wire Mzzow6, Tzzow6, A00pw6, H00pw6, O00pw6, V00pw6, C10pw6, J10pw6, Q10pw6, X10pw6;
wire E20pw6, L20pw6, S20pw6, Z20pw6, G30pw6, N30pw6, U30pw6, B40pw6, I40pw6, P40pw6;
wire W40pw6, D50pw6, K50pw6, R50pw6, Y50pw6, F60pw6, M60pw6, T60pw6, A70pw6, H70pw6;
wire O70pw6, V70pw6, C80pw6, J80pw6, Q80pw6, X80pw6, E90pw6, L90pw6, S90pw6, Z90pw6;
wire Ga0pw6, Na0pw6, Ua0pw6, Bb0pw6, Ib0pw6, Pb0pw6, Wb0pw6, Dc0pw6, Kc0pw6, Rc0pw6;
wire Yc0pw6, Fd0pw6, Md0pw6, Td0pw6, Ae0pw6, He0pw6, Oe0pw6, Ve0pw6, Cf0pw6, Jf0pw6;
wire Qf0pw6, Xf0pw6, Eg0pw6, Lg0pw6, Sg0pw6, Zg0pw6, Gh0pw6, Nh0pw6, Uh0pw6, Bi0pw6;
wire Ii0pw6, Pi0pw6, Wi0pw6, Dj0pw6, Kj0pw6, Rj0pw6, Yj0pw6, Fk0pw6, Mk0pw6, Tk0pw6;
wire Al0pw6, Hl0pw6, Ol0pw6, Vl0pw6, Cm0pw6, Jm0pw6, Qm0pw6, Xm0pw6, En0pw6, Ln0pw6;
wire Sn0pw6, Zn0pw6, Go0pw6, No0pw6, Uo0pw6, Bp0pw6, Ip0pw6, Pp0pw6, Wp0pw6, Dq0pw6;
wire Kq0pw6, Rq0pw6, Yq0pw6, Fr0pw6, Mr0pw6, Tr0pw6, As0pw6, Hs0pw6, Os0pw6, Vs0pw6;
wire Ct0pw6, Jt0pw6, Qt0pw6, Xt0pw6, Eu0pw6, Lu0pw6, Su0pw6, Zu0pw6, Gv0pw6, Nv0pw6;
wire Uv0pw6, Bw0pw6, Iw0pw6, Pw0pw6, Ww0pw6, Dx0pw6, Kx0pw6, Rx0pw6, Yx0pw6, Fy0pw6;
wire My0pw6, Ty0pw6, Az0pw6, Hz0pw6, Oz0pw6, Vz0pw6, C01pw6, J01pw6, Q01pw6, X01pw6;
wire E11pw6, L11pw6, S11pw6, Z11pw6, G21pw6, N21pw6, U21pw6, B31pw6, I31pw6, P31pw6;
wire W31pw6, D41pw6, K41pw6, R41pw6, Y41pw6, F51pw6, M51pw6, T51pw6, A61pw6, H61pw6;
wire O61pw6, V61pw6, C71pw6, J71pw6, Q71pw6, X71pw6, E81pw6, L81pw6, S81pw6, Z81pw6;
wire G91pw6, N91pw6, U91pw6, Ba1pw6, Ia1pw6, Pa1pw6, Wa1pw6, Db1pw6, Kb1pw6, Rb1pw6;
wire Yb1pw6, Fc1pw6, Mc1pw6, Tc1pw6, Ad1pw6, Hd1pw6, Od1pw6, Vd1pw6, Ce1pw6, Je1pw6;
wire Qe1pw6, Xe1pw6, Ef1pw6, Lf1pw6, Sf1pw6, Zf1pw6, Gg1pw6, Ng1pw6, Ug1pw6, Bh1pw6;
wire Ih1pw6, Ph1pw6, Wh1pw6, Di1pw6, Ki1pw6, Ri1pw6, Yi1pw6, Fj1pw6, Mj1pw6, Tj1pw6;
wire Ak1pw6, Hk1pw6, Ok1pw6, Vk1pw6, Cl1pw6, Jl1pw6, Ql1pw6, Xl1pw6, Em1pw6, Lm1pw6;
wire Sm1pw6, Zm1pw6, Gn1pw6, Nn1pw6, Un1pw6, Bo1pw6, Io1pw6, Po1pw6, Wo1pw6, Dp1pw6;
wire Kp1pw6, Rp1pw6, Yp1pw6, Fq1pw6, Mq1pw6, Tq1pw6, Ar1pw6, Hr1pw6, Or1pw6, Vr1pw6;
wire Cs1pw6, Js1pw6, Qs1pw6, Xs1pw6, Et1pw6, Lt1pw6, St1pw6, Zt1pw6, Gu1pw6, Nu1pw6;
wire Uu1pw6, Bv1pw6, Iv1pw6, Pv1pw6, Wv1pw6, Dw1pw6, Kw1pw6, Rw1pw6, Yw1pw6, Fx1pw6;
wire Mx1pw6, Tx1pw6, Ay1pw6, Hy1pw6, Oy1pw6, Vy1pw6, Cz1pw6, Jz1pw6, Qz1pw6, Xz1pw6;
wire E02pw6, L02pw6, S02pw6, Z02pw6, G12pw6, N12pw6, U12pw6, B22pw6, I22pw6, P22pw6;
wire W22pw6, D32pw6, K32pw6, R32pw6, Y32pw6, F42pw6, M42pw6, T42pw6, A52pw6, H52pw6;
wire O52pw6, V52pw6, C62pw6, J62pw6, Q62pw6, X62pw6, E72pw6, L72pw6, S72pw6, Z72pw6;
wire G82pw6, N82pw6, U82pw6, B92pw6, I92pw6, P92pw6, W92pw6, Da2pw6, Ka2pw6, Ra2pw6;
wire Ya2pw6, Fb2pw6, Mb2pw6, Tb2pw6, Ac2pw6, Hc2pw6, Oc2pw6, Vc2pw6, Cd2pw6, Jd2pw6;
wire Qd2pw6, Xd2pw6, Ee2pw6, Le2pw6, Se2pw6, Ze2pw6, Gf2pw6, Nf2pw6, Uf2pw6, Bg2pw6;
wire Ig2pw6, Pg2pw6, Wg2pw6, Dh2pw6, Kh2pw6, Rh2pw6, Yh2pw6, Fi2pw6, Mi2pw6, Ti2pw6;
wire Aj2pw6, Hj2pw6, Oj2pw6, Vj2pw6, Ck2pw6, Jk2pw6, Qk2pw6, Xk2pw6, El2pw6, Ll2pw6;
wire Sl2pw6, Zl2pw6, Gm2pw6, Nm2pw6, Um2pw6, Bn2pw6, In2pw6, Pn2pw6, Wn2pw6, Do2pw6;
wire Ko2pw6, Ro2pw6, Yo2pw6, Fp2pw6, Mp2pw6, Tp2pw6, Aq2pw6, Hq2pw6, Oq2pw6, Vq2pw6;
wire Cr2pw6, Jr2pw6, Qr2pw6, Xr2pw6, Es2pw6, Ls2pw6, Ss2pw6, Zs2pw6, Gt2pw6, Nt2pw6;
wire Ut2pw6, Bu2pw6, Iu2pw6, Pu2pw6, Wu2pw6, Dv2pw6, Kv2pw6, Rv2pw6, Yv2pw6, Fw2pw6;
wire Mw2pw6, Tw2pw6, Ax2pw6, Hx2pw6, Ox2pw6, Vx2pw6, Cy2pw6, Jy2pw6, Qy2pw6, Xy2pw6;
wire Ez2pw6, Lz2pw6, Sz2pw6, Zz2pw6, G03pw6, N03pw6, U03pw6, B13pw6, I13pw6, P13pw6;
wire W13pw6, D23pw6, K23pw6, R23pw6, Y23pw6, F33pw6, M33pw6, T33pw6, A43pw6, H43pw6;
wire O43pw6, V43pw6, C53pw6, J53pw6, Q53pw6, X53pw6, E63pw6, L63pw6, S63pw6, Z63pw6;
wire G73pw6, N73pw6, U73pw6, B83pw6, I83pw6, P83pw6, W83pw6, D93pw6, K93pw6, R93pw6;
wire Y93pw6, Fa3pw6, Ma3pw6, Ta3pw6, Ab3pw6, Hb3pw6, Ob3pw6, Vb3pw6, Cc3pw6, Jc3pw6;
wire Qc3pw6, Xc3pw6, Ed3pw6, Ld3pw6, Sd3pw6, Zd3pw6, Ge3pw6, Ne3pw6, Ue3pw6, Bf3pw6;
wire If3pw6, Pf3pw6, Wf3pw6, Dg3pw6, Kg3pw6, Rg3pw6, Yg3pw6, Fh3pw6, Mh3pw6, Th3pw6;
wire Ai3pw6, Hi3pw6, Oi3pw6, Vi3pw6, Cj3pw6, Jj3pw6, Qj3pw6, Xj3pw6, Ek3pw6, Lk3pw6;
wire Sk3pw6, Zk3pw6, Gl3pw6, Nl3pw6, Ul3pw6, Bm3pw6, Im3pw6, Pm3pw6, Wm3pw6, Dn3pw6;
wire Kn3pw6, Rn3pw6, Yn3pw6, Fo3pw6, Mo3pw6, To3pw6, Ap3pw6, Hp3pw6, Op3pw6, Vp3pw6;
wire Cq3pw6, Jq3pw6, Qq3pw6, Xq3pw6, Er3pw6, Lr3pw6, Sr3pw6, Zr3pw6, Gs3pw6, Ns3pw6;
wire Us3pw6, Bt3pw6, It3pw6, Pt3pw6, Wt3pw6, Du3pw6, Ku3pw6, Ru3pw6, Yu3pw6, Fv3pw6;
wire Mv3pw6, Tv3pw6, Aw3pw6, Hw3pw6, Ow3pw6, Vw3pw6, Cx3pw6, Jx3pw6, Qx3pw6, Xx3pw6;
wire Ey3pw6, Ly3pw6, Sy3pw6, Zy3pw6, Gz3pw6, Nz3pw6, Uz3pw6, B04pw6, I04pw6, P04pw6;
wire W04pw6, D14pw6, K14pw6, R14pw6, Y14pw6, F24pw6, M24pw6, T24pw6, A34pw6, H34pw6;
wire O34pw6, V34pw6, C44pw6, J44pw6, Q44pw6, X44pw6, E54pw6, L54pw6, S54pw6, Z54pw6;
wire G64pw6, N64pw6, U64pw6, B74pw6, I74pw6, P74pw6, W74pw6, D84pw6, K84pw6, R84pw6;
wire Y84pw6, F94pw6, M94pw6, T94pw6, Aa4pw6, Ha4pw6, Oa4pw6, Va4pw6, Cb4pw6, Jb4pw6;
wire Qb4pw6, Xb4pw6, Ec4pw6, Lc4pw6, Sc4pw6, Zc4pw6, Gd4pw6, Nd4pw6, Ud4pw6, Be4pw6;
wire Ie4pw6, Pe4pw6, We4pw6, Df4pw6, Kf4pw6, Rf4pw6, Yf4pw6, Fg4pw6, Mg4pw6, Tg4pw6;
wire Ah4pw6, Hh4pw6, Oh4pw6, Vh4pw6, Ci4pw6, Ji4pw6, Qi4pw6, Xi4pw6, Ej4pw6, Lj4pw6;
wire Sj4pw6, Zj4pw6, Gk4pw6, Nk4pw6, Uk4pw6, Bl4pw6, Il4pw6, Pl4pw6, Wl4pw6, Dm4pw6;
wire Km4pw6, Rm4pw6, Ym4pw6, Fn4pw6, Mn4pw6, Tn4pw6, Ao4pw6, Ho4pw6, Oo4pw6, Vo4pw6;
wire Cp4pw6, Jp4pw6, Qp4pw6, Xp4pw6, Eq4pw6, Lq4pw6, Sq4pw6, Zq4pw6, Gr4pw6, Nr4pw6;
wire Ur4pw6, Bs4pw6, Is4pw6, Ps4pw6, Ws4pw6, Dt4pw6, Kt4pw6, Rt4pw6, Yt4pw6, Fu4pw6;
wire Mu4pw6, Tu4pw6, Av4pw6, Hv4pw6, Ov4pw6, Vv4pw6, Cw4pw6, Jw4pw6, Qw4pw6, Xw4pw6;
wire Ex4pw6, Lx4pw6, Sx4pw6, Zx4pw6, Gy4pw6, Ny4pw6, Uy4pw6, Bz4pw6, Iz4pw6, Pz4pw6;
wire Wz4pw6, D05pw6, K05pw6, R05pw6, Y05pw6, F15pw6, M15pw6, T15pw6, A25pw6, H25pw6;
wire O25pw6, V25pw6, C35pw6, J35pw6, Q35pw6, X35pw6, E45pw6, L45pw6, S45pw6, Z45pw6;
wire G55pw6, N55pw6, U55pw6, B65pw6, I65pw6, P65pw6, W65pw6, D75pw6, K75pw6, R75pw6;
wire Y75pw6, F85pw6, M85pw6, T85pw6, A95pw6, H95pw6, O95pw6, V95pw6, Ca5pw6, Ja5pw6;
wire Qa5pw6, Xa5pw6, Eb5pw6, Lb5pw6, Sb5pw6, Zb5pw6, Gc5pw6, Nc5pw6, Uc5pw6, Bd5pw6;
wire Id5pw6, Pd5pw6, Wd5pw6, De5pw6, Ke5pw6, Re5pw6, Ye5pw6, Ff5pw6, Mf5pw6, Tf5pw6;
wire Ag5pw6, Hg5pw6, Og5pw6, Vg5pw6, Ch5pw6, Jh5pw6, Qh5pw6, Xh5pw6, Ei5pw6, Li5pw6;
wire Si5pw6, Zi5pw6, Gj5pw6, Nj5pw6, Uj5pw6, Bk5pw6, Ik5pw6, Pk5pw6, Wk5pw6, Dl5pw6;
wire Kl5pw6, Rl5pw6, Yl5pw6, Fm5pw6, Mm5pw6, Tm5pw6, An5pw6, Hn5pw6, On5pw6, Vn5pw6;
wire Co5pw6, Jo5pw6, Qo5pw6, Xo5pw6, Ep5pw6, Lp5pw6, Sp5pw6, Zp5pw6, Gq5pw6, Nq5pw6;
wire Uq5pw6, Br5pw6, Ir5pw6, Pr5pw6, Wr5pw6, Ds5pw6, Ks5pw6, Rs5pw6, Ys5pw6, Ft5pw6;
wire Mt5pw6, Tt5pw6, Au5pw6, Hu5pw6, Ou5pw6, Vu5pw6, Cv5pw6, Jv5pw6, Qv5pw6, Xv5pw6;
wire Ew5pw6, Lw5pw6, Sw5pw6, Zw5pw6, Gx5pw6, Nx5pw6, Ux5pw6, By5pw6, Iy5pw6, Py5pw6;
wire Wy5pw6, Dz5pw6, Kz5pw6, Rz5pw6, Yz5pw6, F06pw6, M06pw6, T06pw6, A16pw6, H16pw6;
wire O16pw6, V16pw6, C26pw6, J26pw6, Q26pw6, X26pw6, E36pw6, L36pw6, S36pw6, Z36pw6;
wire G46pw6, N46pw6, U46pw6, B56pw6, I56pw6, P56pw6, W56pw6, D66pw6, K66pw6, R66pw6;
wire Y66pw6, F76pw6, M76pw6, T76pw6, A86pw6, H86pw6, O86pw6, V86pw6, C96pw6, J96pw6;
wire Q96pw6, X96pw6, Ea6pw6, La6pw6, Sa6pw6, Za6pw6, Gb6pw6, Nb6pw6, Ub6pw6, Bc6pw6;
wire Ic6pw6, Pc6pw6, Wc6pw6, Dd6pw6, Kd6pw6, Rd6pw6, Yd6pw6, Fe6pw6, Me6pw6, Te6pw6;
wire Af6pw6, Hf6pw6, Of6pw6, Vf6pw6, Cg6pw6, Jg6pw6, Qg6pw6, Xg6pw6, Eh6pw6, Lh6pw6;
wire Sh6pw6, Zh6pw6, Gi6pw6, Ni6pw6, Ui6pw6, Bj6pw6, Ij6pw6, Pj6pw6, Wj6pw6, Dk6pw6;
wire Kk6pw6, Rk6pw6, Yk6pw6, Fl6pw6, Ml6pw6, Tl6pw6, Am6pw6, Hm6pw6, Om6pw6, Vm6pw6;
wire Cn6pw6, Jn6pw6, Qn6pw6, Xn6pw6, Eo6pw6, Lo6pw6, So6pw6, Zo6pw6, Gp6pw6, Np6pw6;
wire Up6pw6, Bq6pw6, Iq6pw6, Pq6pw6, Wq6pw6, Dr6pw6, Kr6pw6, Rr6pw6, Yr6pw6, Fs6pw6;
wire Ms6pw6, Ts6pw6, At6pw6, Ht6pw6, Ot6pw6, Vt6pw6, Cu6pw6, Ju6pw6, Qu6pw6, Xu6pw6;
wire Ev6pw6, Lv6pw6, Sv6pw6, Zv6pw6, Gw6pw6, Nw6pw6, Uw6pw6, Bx6pw6, Ix6pw6, Px6pw6;
wire Wx6pw6, Dy6pw6, Ky6pw6, Ry6pw6, Yy6pw6, Fz6pw6, Mz6pw6, Tz6pw6, A07pw6, H07pw6;
wire O07pw6, V07pw6, C17pw6, J17pw6, Q17pw6, X17pw6, E27pw6, L27pw6, S27pw6, Z27pw6;
wire G37pw6, N37pw6, U37pw6, B47pw6, I47pw6, P47pw6, W47pw6, D57pw6, K57pw6, R57pw6;
wire Y57pw6, F67pw6, M67pw6, T67pw6, A77pw6, H77pw6, O77pw6, V77pw6, C87pw6, J87pw6;
wire Q87pw6, X87pw6, E97pw6, L97pw6, S97pw6, Z97pw6, Ga7pw6, Na7pw6, Ua7pw6, Bb7pw6;
wire Ib7pw6, Pb7pw6, Wb7pw6, Dc7pw6, Kc7pw6, Rc7pw6, Yc7pw6, Fd7pw6, Md7pw6, Td7pw6;
wire Ae7pw6, He7pw6, Oe7pw6, Ve7pw6, Cf7pw6, Jf7pw6, Qf7pw6, Xf7pw6, Eg7pw6, Lg7pw6;
wire Sg7pw6, Zg7pw6, Gh7pw6, Nh7pw6, Uh7pw6, Bi7pw6, Ii7pw6, Pi7pw6, Wi7pw6, Dj7pw6;
wire Kj7pw6, Rj7pw6, Yj7pw6, Fk7pw6, Mk7pw6, Tk7pw6, Al7pw6, Hl7pw6, Ol7pw6, Vl7pw6;
wire Cm7pw6, Jm7pw6, Qm7pw6, Xm7pw6, En7pw6, Ln7pw6, Sn7pw6, Zn7pw6, Go7pw6, No7pw6;
wire Uo7pw6, Bp7pw6, Ip7pw6, Pp7pw6, Wp7pw6, Dq7pw6, Kq7pw6, Rq7pw6, Yq7pw6, Fr7pw6;
wire Mr7pw6, Tr7pw6, As7pw6, Hs7pw6, Os7pw6, Vs7pw6, Ct7pw6, Jt7pw6, Qt7pw6, Xt7pw6;
wire Eu7pw6, Lu7pw6, Su7pw6, Zu7pw6, Gv7pw6, Nv7pw6, Uv7pw6, Bw7pw6, Iw7pw6, Pw7pw6;
wire Ww7pw6, Dx7pw6, Kx7pw6, Rx7pw6, Yx7pw6, Fy7pw6, My7pw6, Ty7pw6, Az7pw6, Hz7pw6;
wire Oz7pw6, Vz7pw6, C08pw6, J08pw6, Q08pw6, X08pw6, E18pw6, L18pw6, S18pw6, Z18pw6;
wire G28pw6, N28pw6, U28pw6, B38pw6, I38pw6, P38pw6, W38pw6, D48pw6, K48pw6, R48pw6;
wire Y48pw6, F58pw6, M58pw6, T58pw6, A68pw6, H68pw6, O68pw6, V68pw6, C78pw6, J78pw6;
wire Q78pw6, X78pw6, E88pw6, L88pw6, S88pw6, Z88pw6, G98pw6, N98pw6, U98pw6, Ba8pw6;
wire Ia8pw6, Pa8pw6, Wa8pw6, Db8pw6, Kb8pw6, Rb8pw6, Yb8pw6, Fc8pw6, Mc8pw6, Tc8pw6;
wire Ad8pw6, Hd8pw6, Od8pw6, Vd8pw6, Ce8pw6, Je8pw6, Qe8pw6, Xe8pw6, Ef8pw6, Lf8pw6;
wire Sf8pw6, Zf8pw6, Gg8pw6, Ng8pw6, Ug8pw6, Bh8pw6, Ih8pw6, Ph8pw6, Wh8pw6, Di8pw6;
wire Ki8pw6, Ri8pw6, Yi8pw6, Fj8pw6, Mj8pw6, Tj8pw6, Ak8pw6, Hk8pw6, Ok8pw6, Vk8pw6;
wire Cl8pw6, Jl8pw6, Ql8pw6, Xl8pw6, Em8pw6, Lm8pw6, Sm8pw6, Zm8pw6, Gn8pw6, Nn8pw6;
wire Un8pw6, Bo8pw6, Io8pw6, Po8pw6, Wo8pw6, Dp8pw6, Kp8pw6, Rp8pw6, Yp8pw6, Fq8pw6;
wire Mq8pw6, Tq8pw6, Ar8pw6, Hr8pw6, Or8pw6, Vr8pw6, Cs8pw6, Js8pw6, Qs8pw6, Xs8pw6;
wire Et8pw6, Lt8pw6, St8pw6, Zt8pw6, Gu8pw6, Nu8pw6, Uu8pw6, Bv8pw6, Iv8pw6, Pv8pw6;
wire Wv8pw6, Dw8pw6, Kw8pw6, Rw8pw6, Yw8pw6, Fx8pw6, Mx8pw6, Tx8pw6, Ay8pw6, Hy8pw6;
wire Oy8pw6, Vy8pw6, Cz8pw6, Jz8pw6, Qz8pw6, Xz8pw6, E09pw6, L09pw6, S09pw6, Z09pw6;
wire G19pw6, N19pw6, U19pw6, B29pw6, I29pw6, P29pw6, W29pw6, D39pw6, K39pw6, R39pw6;
wire Y39pw6, F49pw6, M49pw6, T49pw6, A59pw6, H59pw6, O59pw6, V59pw6, C69pw6, J69pw6;
wire Q69pw6, X69pw6, E79pw6, L79pw6, S79pw6, Z79pw6, G89pw6, N89pw6, U89pw6, B99pw6;
wire I99pw6, P99pw6, W99pw6, Da9pw6, Ka9pw6, Ra9pw6, Ya9pw6, Fb9pw6, Mb9pw6, Tb9pw6;
wire Ac9pw6, Hc9pw6, Oc9pw6, Vc9pw6, Cd9pw6, Jd9pw6, Qd9pw6, Xd9pw6, Ee9pw6, Le9pw6;
wire Se9pw6, Ze9pw6, Gf9pw6, Nf9pw6, Uf9pw6, Bg9pw6, Ig9pw6, Pg9pw6, Wg9pw6, Dh9pw6;
wire Kh9pw6, Rh9pw6, Yh9pw6, Fi9pw6, Mi9pw6, Ti9pw6, Aj9pw6, Hj9pw6, Oj9pw6, Vj9pw6;
wire Ck9pw6, Jk9pw6, Qk9pw6, Xk9pw6, El9pw6, Ll9pw6, Sl9pw6, Zl9pw6, Gm9pw6, Nm9pw6;
wire Um9pw6, Bn9pw6, In9pw6, Pn9pw6, Wn9pw6, Do9pw6, Ko9pw6, Ro9pw6, Yo9pw6, Fp9pw6;
wire Mp9pw6, Tp9pw6, Aq9pw6, Hq9pw6, Oq9pw6, Vq9pw6, Cr9pw6, Jr9pw6, Qr9pw6, Xr9pw6;
wire Es9pw6, Ls9pw6, Ss9pw6, Zs9pw6, Gt9pw6, Nt9pw6, Ut9pw6, Bu9pw6, Iu9pw6, Pu9pw6;
wire Wu9pw6, Dv9pw6, Kv9pw6, Rv9pw6, Yv9pw6, Fw9pw6, Mw9pw6, Tw9pw6, Ax9pw6, Hx9pw6;
wire Ox9pw6, Vx9pw6, Cy9pw6, Jy9pw6, Qy9pw6, Xy9pw6, Ez9pw6, Lz9pw6, Sz9pw6, Zz9pw6;
wire G0apw6, N0apw6, U0apw6, B1apw6, I1apw6, P1apw6, W1apw6, D2apw6, K2apw6, R2apw6;
wire Y2apw6, F3apw6, M3apw6, T3apw6, A4apw6, H4apw6, O4apw6, V4apw6, C5apw6, J5apw6;
wire Q5apw6, X5apw6, E6apw6, L6apw6, S6apw6, Z6apw6, G7apw6, N7apw6, U7apw6, B8apw6;
wire I8apw6, P8apw6, W8apw6, D9apw6, K9apw6, R9apw6, Y9apw6, Faapw6, Maapw6, Taapw6;
wire Abapw6, Hbapw6, Obapw6, Vbapw6, Ccapw6, Jcapw6, Qcapw6, Xcapw6, Edapw6, Ldapw6;
wire Sdapw6, Zdapw6, Geapw6, Neapw6, Ueapw6, Bfapw6, Ifapw6, Pfapw6, Wfapw6, Dgapw6;
wire Kgapw6, Rgapw6, Ygapw6, Fhapw6, Mhapw6, Thapw6, Aiapw6, Hiapw6, Oiapw6, Viapw6;
wire Cjapw6, Jjapw6, Qjapw6, Xjapw6, Ekapw6, Lkapw6, Skapw6, Zkapw6, Glapw6, Nlapw6;
wire Ulapw6, Bmapw6, Imapw6, Pmapw6, Wmapw6, Dnapw6, Knapw6, Rnapw6, Ynapw6, Foapw6;
wire Moapw6, Toapw6, Apapw6, Hpapw6, Opapw6, Vpapw6, Cqapw6, Jqapw6, Qqapw6, Xqapw6;
wire Erapw6, Lrapw6, Srapw6, Zrapw6, Gsapw6, Nsapw6, Usapw6, Btapw6, Itapw6, Ptapw6;
wire Wtapw6, Duapw6, Kuapw6, Ruapw6, Yuapw6, Fvapw6, Mvapw6, Tvapw6, Awapw6, Hwapw6;
wire Owapw6, Vwapw6, Cxapw6, Jxapw6, Qxapw6, Xxapw6, Eyapw6, Lyapw6, Syapw6, Zyapw6;
wire Gzapw6, Nzapw6, Uzapw6, B0bpw6, I0bpw6, P0bpw6, W0bpw6, D1bpw6, K1bpw6, R1bpw6;
wire Y1bpw6, F2bpw6, M2bpw6, T2bpw6, A3bpw6, H3bpw6, O3bpw6, V3bpw6, C4bpw6, J4bpw6;
wire Q4bpw6, X4bpw6, E5bpw6, L5bpw6, S5bpw6, Z5bpw6, G6bpw6, N6bpw6, U6bpw6, B7bpw6;
wire I7bpw6, P7bpw6, W7bpw6, D8bpw6, K8bpw6, R8bpw6, Y8bpw6, F9bpw6, M9bpw6, T9bpw6;
wire Aabpw6, Habpw6, Oabpw6, Vabpw6, Cbbpw6, Jbbpw6, Qbbpw6, Xbbpw6, Ecbpw6, Lcbpw6;
wire Scbpw6, Zcbpw6, Gdbpw6, Ndbpw6, Udbpw6, Bebpw6, Iebpw6, Pebpw6, Webpw6, Dfbpw6;
wire Kfbpw6, Rfbpw6, Yfbpw6, Fgbpw6, Mgbpw6, Tgbpw6, Ahbpw6, Hhbpw6, Ohbpw6, Vhbpw6;
wire Cibpw6, Jibpw6, Qibpw6, Xibpw6, Ejbpw6, Ljbpw6, Sjbpw6, Zjbpw6, Gkbpw6, Nkbpw6;
wire Ukbpw6, Blbpw6, Ilbpw6, Plbpw6, Wlbpw6, Dmbpw6, Kmbpw6, Rmbpw6, Ymbpw6, Fnbpw6;
wire Mnbpw6, Tnbpw6, Aobpw6, Hobpw6, Oobpw6, Vobpw6, Cpbpw6, Jpbpw6, Qpbpw6, Xpbpw6;
wire Eqbpw6, Lqbpw6, Sqbpw6, Zqbpw6, Grbpw6, Nrbpw6, Urbpw6, Bsbpw6, Isbpw6, Psbpw6;
wire Wsbpw6, Dtbpw6, Ktbpw6, Rtbpw6, Ytbpw6, Fubpw6, Mubpw6, Tubpw6, Avbpw6, Hvbpw6;
wire Ovbpw6, Vvbpw6, Cwbpw6, Jwbpw6, Qwbpw6, Xwbpw6, Exbpw6, Lxbpw6, Sxbpw6, Zxbpw6;
wire Gybpw6, Nybpw6, Uybpw6, Bzbpw6, Izbpw6, Pzbpw6, Wzbpw6, D0cpw6, K0cpw6, R0cpw6;
wire Y0cpw6, F1cpw6, M1cpw6, T1cpw6, A2cpw6, H2cpw6, O2cpw6, V2cpw6, C3cpw6, J3cpw6;
wire Q3cpw6, X3cpw6, E4cpw6, L4cpw6, S4cpw6, Z4cpw6, G5cpw6, N5cpw6, U5cpw6, B6cpw6;
wire I6cpw6, P6cpw6, W6cpw6, D7cpw6, K7cpw6, R7cpw6, Y7cpw6, F8cpw6, M8cpw6, T8cpw6;
wire A9cpw6, H9cpw6, O9cpw6, V9cpw6, Cacpw6, Jacpw6, Qacpw6, Xacpw6, Ebcpw6, Lbcpw6;
wire Sbcpw6, Zbcpw6, Gccpw6, Nccpw6, Uccpw6, Bdcpw6, Idcpw6, Pdcpw6, Wdcpw6, Decpw6;
wire Kecpw6, Recpw6, Yecpw6, Ffcpw6, Mfcpw6, Tfcpw6, Agcpw6, Hgcpw6, Ogcpw6, Vgcpw6;
wire Chcpw6, Jhcpw6, Qhcpw6, Xhcpw6, Eicpw6, Licpw6, Sicpw6, Zicpw6, Gjcpw6, Njcpw6;
wire Ujcpw6, Bkcpw6, Ikcpw6, Pkcpw6, Wkcpw6, Dlcpw6, Klcpw6, Rlcpw6, Ylcpw6, Fmcpw6;
wire Mmcpw6, Tmcpw6, Ancpw6, Hncpw6, Oncpw6, Vncpw6, Cocpw6, Jocpw6, Qocpw6, Xocpw6;
wire Epcpw6, Lpcpw6, Spcpw6, Zpcpw6, Gqcpw6, Nqcpw6, Uqcpw6, Brcpw6, Ircpw6, Prcpw6;
wire Wrcpw6, Dscpw6, Kscpw6, Rscpw6, Yscpw6, Ftcpw6, Mtcpw6, Ttcpw6, Aucpw6, Hucpw6;
wire Oucpw6, Vucpw6, Cvcpw6, Jvcpw6, Qvcpw6, Xvcpw6, Ewcpw6, Lwcpw6, Swcpw6, Zwcpw6;
wire Gxcpw6, Nxcpw6, Uxcpw6, Bycpw6, Iycpw6, Pycpw6, Wycpw6, Dzcpw6, Kzcpw6, Rzcpw6;
wire Yzcpw6, F0dpw6, M0dpw6, T0dpw6, A1dpw6, H1dpw6, O1dpw6, V1dpw6, C2dpw6, J2dpw6;
wire Q2dpw6, X2dpw6, E3dpw6, L3dpw6, S3dpw6, Z3dpw6, G4dpw6, N4dpw6, U4dpw6, B5dpw6;
wire I5dpw6, P5dpw6, W5dpw6, D6dpw6, K6dpw6, R6dpw6, Y6dpw6, F7dpw6, M7dpw6, T7dpw6;
wire A8dpw6, H8dpw6, O8dpw6, V8dpw6, C9dpw6, J9dpw6, Q9dpw6, X9dpw6, Eadpw6, Ladpw6;
wire Sadpw6, Zadpw6, Gbdpw6, Nbdpw6, Ubdpw6, Bcdpw6, Icdpw6, Pcdpw6, Wcdpw6, Dddpw6;
wire Kddpw6, Rddpw6, Yddpw6, Fedpw6, Medpw6, Tedpw6, Afdpw6, Hfdpw6, Ofdpw6, Vfdpw6;
wire Cgdpw6, Jgdpw6, Qgdpw6, Xgdpw6, Ehdpw6, Lhdpw6, Shdpw6, Zhdpw6, Gidpw6, Nidpw6;
wire Uidpw6, Bjdpw6, Ijdpw6, Pjdpw6, Wjdpw6, Dkdpw6, Kkdpw6, Rkdpw6, Ykdpw6, Fldpw6;
wire Mldpw6, Tldpw6, Amdpw6, Hmdpw6, Omdpw6, Vmdpw6, Cndpw6, Jndpw6, Qndpw6, Xndpw6;
wire Eodpw6, Lodpw6, Sodpw6, Zodpw6, Gpdpw6, Npdpw6, Updpw6, Bqdpw6, Iqdpw6, Pqdpw6;
wire Wqdpw6, Drdpw6, Krdpw6, Rrdpw6, Yrdpw6, Fsdpw6, Msdpw6, Tsdpw6, Atdpw6, Htdpw6;
wire Otdpw6, Vtdpw6, Cudpw6, Judpw6, Qudpw6, Xudpw6, Evdpw6, Lvdpw6, Svdpw6, Zvdpw6;
wire Gwdpw6, Nwdpw6, Uwdpw6, Bxdpw6, Ixdpw6, Pxdpw6, Wxdpw6, Dydpw6, Kydpw6, Rydpw6;
wire Yydpw6, Fzdpw6, Mzdpw6, Tzdpw6, A0epw6, H0epw6, O0epw6, V0epw6, C1epw6, J1epw6;
wire Q1epw6, X1epw6, E2epw6, L2epw6, S2epw6, Z2epw6, G3epw6, N3epw6, U3epw6, B4epw6;
wire I4epw6, P4epw6, W4epw6, D5epw6, K5epw6, H6epw6, E7epw6, B8epw6, Y8epw6, V9epw6;
wire Saepw6, Pbepw6, Mcepw6, Jdepw6, Heepw6, Ffepw6, Dgepw6, Bhepw6, Zhepw6, Xiepw6;
wire Vjepw6, Tkepw6, Rlepw6, Pmepw6, Nnepw6, Loepw6, Jpepw6, Hqepw6, Frepw6, Dsepw6;
wire Btepw6, Ztepw6, Xuepw6, Vvepw6, Twepw6, Rxepw6, Pyepw6, Nzepw6, L0fpw6, J1fpw6;
wire [3:0] H2fpw6;
wire [3:0] X3fpw6;
wire [30:2] N5fpw6;
wire [15:0] D7fpw6;
wire [11:0] S8fpw6;
wire [31:0] Eafpw6;
wire [30:0] Qbfpw6;
wire [31:0] Idfpw6;
wire [31:0] Affpw6;
wire [31:0] Tgfpw6;
wire [31:0] Mifpw6;
wire [31:0] Fkfpw6;
wire [8:1] Xlfpw6;
wire [7:0] Vnfpw6;
wire [16:0] Ppfpw6;
wire [16:0] Hrfpw6;
wire [30:0] Zsfpw6;
wire [1:0] Sufpw6;
wire [1:0] Iwfpw6;
wire [7:0] Cyfpw6;
wire [23:0] Tzfpw6;
wire [1:0] L1gpw6;
wire [1:0] B3gpw6;
wire [63:0] R4gpw6;
wire [23:0] L6gpw6;
wire [1:0] H8gpw6;
wire [23:0] Bagpw6;
wire [31:0] Vbgpw6;
wire [31:0] Odgpw6;
wire [4:0] Jfgpw6;
wire [4:0] Dhgpw6;
wire [28:27] Ligpw6;
wire [28:27] Akgpw6;
wire [28:27] Plgpw6;
wire [28:27] Engpw6;
wire [28:2] Togpw6;
wire [28:2] Gqgpw6;
wire [28:2] Trgpw6;
wire [28:2] Gtgpw6;
wire [13:0] Tugpw6;
wire [2:0] Lwgpw6;
wire [4:0] Aygpw6;
wire [1:0] Pzgpw6;
wire [31:2] E1hpw6;
wire [2:0] R2hpw6;
wire [4:0] G4hpw6;
wire [1:0] V5hpw6;
wire [31:2] K7hpw6;
wire [6:0] X8hpw6;
wire [30:0] Iahpw6;
wire [30:26] Zbhpw6;
wire [3:0] Mdhpw6;
wire [6:0] Zehpw6;
wire [5:0] Ighpw6;
wire [31:0] Shhpw6;
wire [3:0] Cjhpw6;
wire [1:0] Pkhpw6;
wire [9:0] Gmhpw6;
wire [3:0] Tnhpw6;
wire [2:1] Aphpw6;
wire [1:0] Sqhpw6;
wire [31:4] Jshpw6;
wire [31:0] Uthpw6;
reg Evhpw6, Hwhpw6, Kxhpw6, Nyhpw6, T0ipw6, A3ipw6, A5ipw6, W6ipw6, M8ipw6, Qaipw6;
reg Tcipw6, Weipw6, Wgipw6, Xiipw6, Wkipw6, Vmipw6, Uoipw6, Uqipw6, Usipw6, Vuipw6;
reg Uwipw6, Tyipw6, V0jpw6, X2jpw6, X4jpw6, X6jpw6, Z8jpw6, Bbjpw6, Bdjpw6, Bfjpw6;
reg Vgjpw6, Qijpw6, Kkjpw6, Kmjpw6, Kojpw6, Lqjpw6, Isjpw6, Aujpw6, Yvjpw6, Wxjpw6;
reg Vzjpw6, U1kpw6, T3kpw6, S5kpw6, R7kpw6, T9kpw6, Vbkpw6, Rdkpw6, Rfkpw6, Rhkpw6;
reg Tjkpw6, Vlkpw6, Vnkpw6, Vpkpw6, Nrkpw6, Stkpw6, Jvkpw6, Oxkpw6, Pzkpw6, I1lpw6;
reg H3lpw6, L5lpw6, B7lpw6, Y8lpw6, Kalpw6, Bclpw6, Sdlpw6, Jflpw6, Ahlpw6, Rilpw6;
reg Yklpw6, Pmlpw6, Golpw6, Vplpw6, Krlpw6, Zslpw6, Oulpw6, Kwlpw6, Gylpw6, Yzlpw6;
reg O1mpw6, S3mpw6, T5mpw6, S7mpw6, R9mpw6, Qbmpw6, Pdmpw6, Ofmpw6, Qhmpw6, Mjmpw6;
reg Mlmpw6, Mnmpw6, Jpmpw6, Irmpw6, Htmpw6, Gvmpw6, Gxmpw6, Fzmpw6, E1npw6, E3npw6;
reg E5npw6, E7npw6, E9npw6, Ebnpw6, Ednpw6, Efnpw6, Ehnpw6, Ejnpw6, Elnpw6, Fnnpw6;
reg Fpnpw6, Arnpw6, Usnpw6, Uunpw6, Zwnpw6, Qynpw6, I0opw6, D2opw6, T3opw6, X5opw6;
reg Y7opw6, Z9opw6, Xbopw6, Ydopw6, Ufopw6, Shopw6, Rjopw6, Qlopw6, Qnopw6, Qpopw6;
reg Propw6, Otopw6, Ovopw6, Oxopw6, Ozopw6, O1ppw6, O3ppw6, O5ppw6, N7ppw6, N9ppw6;
reg Nbppw6, Mdppw6, Lfppw6, Lhppw6, Ljppw6, Llppw6, Lnppw6, Lpppw6, Lrppw6, Ktppw6;
reg Jvppw6, Ixppw6, Izppw6, I1qpw6, I3qpw6, I5qpw6, I7qpw6, I9qpw6, Ibqpw6, Idqpw6;
reg Nfqpw6, Ehqpw6, Cjqpw6, Xkqpw6, Gnqpw6, Gpqpw6, Nrqpw6, Utqpw6, Xvqpw6, Xxqpw6;
reg Yzqpw6, D2rpw6, I4rpw6, M6rpw6, N8rpw6, Oarpw6, Pcrpw6, Lerpw6, Hgrpw6, Hirpw6;
reg Fkrpw6, Emrpw6, Dorpw6, Cqrpw6, Bsrpw6, Aurpw6, Zvrpw6, Yxrpw6, B0spw6, A2spw6;
reg Z3spw6, Y5spw6, X7spw6, W9spw6, Vbspw6, Xdspw6, Wfspw6, Vhspw6, Ujspw6, Wlspw6;
reg Ynspw6, Ypspw6, Yrspw6, Ytspw6, Yvspw6, Yxspw6, Yzspw6, Z1tpw6, Z3tpw6, Z5tpw6;
reg Z7tpw6, Z9tpw6, Zbtpw6, Zdtpw6, Yftpw6, Xhtpw6, Wjtpw6, Vltpw6, Untpw6, Tptpw6;
reg Vrtpw6, Xttpw6, Xvtpw6, Xxtpw6, Xztpw6, X1upw6, X3upw6, X5upw6, Y7upw6, Y9upw6;
reg Ybupw6, Ydupw6, Yfupw6, Yhupw6, Yjupw6, Amupw6, Coupw6, Equpw6, Asupw6, Ztupw6;
reg Awupw6, Xxupw6, Vzupw6, T1vpw6, R3vpw6, P5vpw6, K7vpw6, F9vpw6, Gbvpw6, Ldvpw6;
reg Cfvpw6, Hhvpw6, Jjvpw6, Jlvpw6, Jnvpw6, Jpvpw6, Jrvpw6, Jtvpw6, Jvvpw6, Dxvpw6;
reg Dzvpw6, C1wpw6, C3wpw6, C5wpw6, C7wpw6, C9wpw6, Cbwpw6, Cdwpw6, Cfwpw6, Chwpw6;
reg Cjwpw6, Hlwpw6, Ymwpw6, Dpwpw6, Sqwpw6, Kswpw6, Puwpw6, Gwwpw6, Lywpw6, N0xpw6;
reg P2xpw6, P4xpw6, P6xpw6, P8xpw6, Paxpw6, Pcxpw6, Pexpw6, Jgxpw6, Iixpw6, Hkxpw6;
reg Hmxpw6, Hoxpw6, Hqxpw6, Hsxpw6, Huxpw6, Gwxpw6, Gyxpw6, L0ypw6, C2ypw6, H4ypw6;
reg W5ypw6, X7ypw6, U9ypw6, Ubypw6, Tdypw6, Sfypw6, Rhypw6, Qjypw6, Plypw6, Onypw6;
reg Npypw6, Jrypw6, Ftypw6, Evypw6, Exypw6, Ezypw6, D1zpw6, C3zpw6, B5zpw6, A7zpw6;
reg Z8zpw6, Zazpw6, Zczpw6, Zezpw6, Zgzpw6, Yizpw6, Ykzpw6, Ymzpw6, Xozpw6, Wqzpw6;
reg Vszpw6, Uuzpw6, Twzpw6, Tyzpw6, T00qw6, T20qw6, T40qw6, T60qw6, T80qw6, Ta0qw6;
reg Tc0qw6, Te0qw6, Tg0qw6, Ti0qw6, Tk0qw6, Tm0qw6, So0qw6, Rq0qw6, Ss0qw6, Tu0qw6;
reg Sw0qw6, Ry0qw6, Q01qw6, P21qw6, O41qw6, N61qw6, M81qw6, Qa1qw6, Gc1qw6, Ke1qw6;
reg Yf1qw6, Mh1qw6, Qj1qw6, Gl1qw6, Kn1qw6, Jp1qw6, Ir1qw6, Ht1qw6, Gv1qw6, Fx1qw6;
reg Ez1qw6, D12qw6, A32qw6, X42qw6, C72qw6, T82qw6, Ra2qw6, Wc2qw6, Le2qw6, Dg2qw6;
reg Uh2qw6, Nj2qw6, Fl2qw6, Kn2qw6, Bp2qw6, Gr2qw6, Bt2qw6, Xu2qw6, Bx2qw6, Ry2qw6;
reg L03qw6, P23qw6, D43qw6, V53qw6, Z73qw6, P93qw6, Tb3qw6, Nd3qw6, Bf3qw6, Pg3qw6;
reg Di3qw6, Vj3qw6, Jl3qw6, Ym3qw6, No3qw6, Cq3qw6, Rr3qw6, Wt3qw6, Nv3qw6, Sx3qw6;
reg Sz3qw6, P14qw6, P34qw6, P54qw6, Gp6ax6, Gr6ax6, Gt6ax6, Gv6ax6, Gx6ax6, Gz6ax6;
reg F17ax6, C37ax6, Z47ax6, Z67ax6, E97ax6, Va7ax6, Ad7ax6, Pe7ax6, Hg7ax6, Li7ax6;
reg Bk7ax6, Fm7ax6, Xn7ax6, Lp7ax6, Nr7ax6, Pt7ax6, Rv7ax6, Sx7ax6, Sz7ax6, S18ax6;
reg S38ax6, S58ax6, S78ax6, S98ax6, Sb8ax6, Sd8ax6, Xf8ax6, Oh8ax6, Fj8ax6, Kl8ax6;
reg Zm8ax6, Ro8ax6, Wq8ax6, Ns8ax6, Su8ax6, Hw8ax6, Zx8ax6, Vz8ax6, R19ax6, N39ax6;
reg J59ax6, G79ax6, D99ax6, Ab9ax6, Xc9ax6, Ue9ax6, Rg9ax6, Oi9ax6, Lk9ax6, Im9ax6;
reg Fo9ax6, Bq9ax6, Xr9ax6, Tt9ax6, Pv9ax6, Lx9ax6, Hz9ax6, D1aax6, Z2aax6, W4aax6;
reg T6aax6, Q8aax6, Naaax6, Kcaax6, Heaax6, Egaax6, Biaax6, Yjaax6, Vlaax6, Rnaax6;
reg Npaax6, Jraax6, Ftaax6, Bvaax6, Xwaax6, Tyaax6, P0bax6, L2bax6, H4bax6, X5bax6;
reg T7bax6, P9bax6, Lbbax6, Hdbax6, Dfbax6, Zgbax6, Vibax6, Rkbax6, Hmbax6, Xnbax6;
reg Opbax6, Krbax6, Htbax6, Evbax6, Bxbax6, Yybax6, V0cax6, S2cax6, P4cax6, M6cax6;
reg J8cax6, Facax6, Bccax6, Xdcax6, Tfcax6, Phcax6, Ljcax6, Hlcax6, Dncax6, Apcax6;
reg Xqcax6, Uscax6, Rucax6, Owcax6, Lycax6, I0dax6, F2dax6, C4dax6, Y5dax6, U7dax6;
reg Q9dax6, Mbdax6, Iddax6, Efdax6, Ahdax6, Widax6, Tkdax6, Qmdax6, Nodax6, Kqdax6;
reg Hsdax6, Eudax6, Bwdax6, Yxdax6, Vzdax6, R1eax6, N3eax6, J5eax6, F7eax6, B9eax6;
reg Xaeax6, Tceax6, Peeax6, Mgeax6, Jieax6, Gkeax6, Dmeax6, Aoeax6, Xpeax6, Ureax6;
reg Rteax6, Oveax6, Kxeax6, Gzeax6, C1fax6, Y2fax6, U4fax6, Q6fax6, M8fax6, Eafax6;
reg Sbfax6, Hdfax6, Vefax6, Zgfax6, Pifax6, Okfax6, Nmfax6, Uofax6, Sqfax6, Qsfax6;
reg Qufax6, Qwfax6, Ryfax6, J0gax6, Q2gax6, N4gax6, K6gax6, H8gax6, Eagax6, Bcgax6;
reg Ydgax6, Nfgax6, Khgax6, Hjgax6, Elgax6, Bngax6, Yogax6, Vqgax6, Ksgax6, Dugax6;
reg Wvgax6, Jxgax6, Vygax6, U0hax6, R2hax6, O4hax6, L6hax6, I8hax6, Fahax6, Cchax6;
reg Zdhax6, Wfhax6, Thhax6, Qjhax6, Nlhax6, Knhax6, Hphax6, Drhax6, Zshax6, Vuhax6;
reg Rwhax6, Nyhax6, J0iax6, G2iax6, F4iax6, E6iax6, E8iax6, Daiax6, Bciax6, Zdiax6;
reg Xfiax6, Thiax6, Ijiax6, Eliax6, Aniax6, Woiax6, Zqiax6, Ysiax6, Xuiax6, Wwiax6;
reg Wyiax6, W0jax6, W2jax6, W4jax6, V6jax6, U8jax6, Tajax6, Tcjax6, Sejax6, Sgjax6;
reg Sijax6, Skjax6, Smjax6, Sojax6, Sqjax6, Ssjax6, Sujax6, Rwjax6, Qyjax6, P0kax6;
reg O2kax6, N4kax6, M6kax6, L8kax6, Kakax6, Jckax6, Iekax6, Lgkax6, Oikax6, Rkkax6;
reg Umkax6, Tokax6, Sqkax6, Rskax6, Qukax6, Pwkax6, Oykax6, N0lax6, M2lax6, L4lax6;
reg L6lax6, I8lax6, Halax6, Eclax6, Delax6, Cglax6, Cilax6, Cklax6, Cmlax6, Bolax6;
reg Aqlax6, Zrlax6, Ytlax6, Xvlax6, Xxlax6, Xzlax6, X1max6, X3max6, W5max6, W7max6;
reg W9max6, Wbmax6, Wdmax6, Wfmax6, Whmax6, Wjmax6, Wlmax6, Wnmax6, Wpmax6, Wrmax6;
reg Vtmax6, Uvmax6, Txmax6, Szmax6, S1nax6, S3nax6, S5nax6, R7nax6, Q9nax6, Pbnax6;
reg Odnax6, Nfnax6, Nhnax6, Njnax6, Nlnax6, Nnnax6, Npnax6, Nrnax6, Ntnax6, Nvnax6;
reg Nxnax6, Nznax6, N1oax6, N3oax6, N5oax6, N7oax6, N9oax6, Mboax6, Ldoax6, Kfoax6;
reg Khoax6, Kjoax6, Kloax6, Jnoax6, Ipoax6, Hroax6, Gtoax6, Fvoax6, Fxoax6, Fzoax6;
reg F1pax6, F3pax6, E5pax6, E7pax6, E9pax6, Ebpax6, Edpax6, Efpax6, Ehpax6, Ejpax6;
reg Elpax6, Enpax6, Eppax6, Erpax6, Dtpax6, Cvpax6, Bxpax6, Azpax6, A1qax6, A3qax6;
reg A5qax6, Z6qax6, Y8qax6, Xaqax6, Wcqax6, Veqax6, Vgqax6, Viqax6, Vkqax6, Vmqax6;
reg Uoqax6, Uqqax6, Usqax6, Uuqax6, Uwqax6, Uyqax6, U0rax6, U2rax6, U4rax6, U6rax6;
reg U8rax6, Uarax6, Tcrax6, Serax6, Rgrax6, Qirax6, Qkrax6, Qmrax6, Qorax6, Pqrax6;
reg Osrax6, Ourax6, Owrax6, Oyrax6, O0sax6, O2sax6, O4sax6, O6sax6, O8sax6, Oasax6;
reg Ocsax6, Oesax6, Ngsax6, Misax6, Lksax6, Kmsax6, Kosax6, Kqsax6, Kssax6, Jusax6;
reg Iwsax6, Hysax6, G0tax6, F2tax6, F4tax6, F6tax6, F8tax6, Fatax6, Ectax6, Eetax6;
reg Egtax6, Eitax6, Ektax6, Emtax6, Eotax6, Eqtax6, Estax6, Eutax6, Ewtax6, Eytax6;
reg D0uax6, C2uax6, B4uax6, B6uax6, B8uax6, Bauax6, Acuax6, Zduax6, Yfuax6, Xhuax6;
reg Wjuax6, Wluax6, Wnuax6, Wpuax6, Wruax6, Vtuax6, Vvuax6, Vxuax6, Vzuax6, V1vax6;
reg V3vax6, V5vax6, V7vax6, V9vax6, Vbvax6, Vdvax6, Vfvax6, Uhvax6, Tjvax6, Slvax6;
reg Rnvax6, Rpvax6, Rrvax6, Rtvax6, Qvvax6, Pxvax6, Ozvax6, N1wax6, M3wax6, M5wax6;
reg M7wax6, M9wax6, Mbwax6, Ldwax6, Lfwax6, Lhwax6, Ljwax6, Llwax6, Lnwax6, Lpwax6;
reg Lrwax6, Ltwax6, Lvwax6, Lxwax6, Lzwax6, K1xax6, J3xax6, I5xax6, J7xax6, L9xax6;
reg Nbxax6, Pdxax6, Rfxax6, Thxax6, Ujxax6, Vlxax6, Wnxax6, Xpxax6, Xrxax6, Wtxax6;
reg Vvxax6, Vxxax6, Vzxax6, V1yax6, U3yax6, T5yax6, S7yax6, R9yax6, Sbyax6, Pdyax6;
reg Mfyax6, Ohyax6, Qjyax6, Slyax6, Unyax6, Wpyax6, Yryax6, Auyax6, Cwyax6, Eyyax6;
reg G0zax6, I2zax6, H4zax6, J6zax6, L8zax6, Nazax6, Pczax6, Rezax6, Tgzax6, Uizax6;
reg Vkzax6, Wmzax6, Xozax6, Yqzax6, Zszax6, Avzax6, Cxzax6, Czzax6, C10bx6, C30bx6;
reg C50bx6, D70bx6, E90bx6, Fb0bx6, Gd0bx6, Hf0bx6, Ih0bx6, Jj0bx6, Kl0bx6, Ln0bx6;
reg Mp0bx6, Nr0bx6, Ot0bx6, Pv0bx6, Qx0bx6, Rz0bx6, S11bx6, U31bx6, W51bx6, Z71bx6;
reg Ca1bx6, Fc1bx6, Ie1bx6, Lg1bx6, Oi1bx6, Rk1bx6, Um1bx6, Xo1bx6, Ar1bx6, Dt1bx6;
reg Gv1bx6, Jx1bx6, Mz1bx6, P12bx6, S32bx6, V52bx6, Y72bx6, Aa2bx6, Cc2bx6, Fe2bx6;
reg Ig2bx6, Li2bx6, Ok2bx6, Rm2bx6, Uo2bx6, Xq2bx6, At2bx6, Dv2bx6, Gx2bx6, Jz2bx6;
reg M13bx6, P33bx6, S53bx6, V73bx6, Y93bx6, Bc3bx6, Ee3bx6, Hg3bx6, Ki3bx6, Mk3bx6;
reg Om3bx6, Qo3bx6, Sq3bx6, Us3bx6, Wu3bx6, Yw3bx6, Az3bx6, C14bx6, E34bx6, G54bx6;
reg I74bx6, K94bx6, Mb4bx6, Od4bx6, Qf4bx6, Sh4bx6, Uj4bx6, Tl4bx6, Sn4bx6, Up4bx6;
reg Wr4bx6, Yt4bx6, Aw4bx6, Cy4bx6, E05bx6, G25bx6, I45bx6, K65bx6, M85bx6, Oa5bx6;
reg Qc5bx6, Pe5bx6, Og5bx6, Ni5bx6, Nk5bx6, Nm5bx6, No5bx6, Nq5bx6, Ms5bx6, Nu5bx6;
reg Mw5bx6, Jy5bx6, J06bx6, F26bx6, D46bx6, D66bx6, D86bx6, Da6bx6, Dc6bx6, De6bx6;
reg Dg6bx6, Di6bx6, Dk6bx6, Dm6bx6, Do6bx6, Dq6bx6, Cs6bx6, Bu6bx6, Gw6bx6, Xx6bx6;
reg C07bx6, C27bx6, C47bx6, C67bx6, C87bx6, Ca7bx6, Cc7bx6, Ce7bx6, Cg7bx6, Ci7bx6;
reg Ck7bx6, Cm7bx6, Co7bx6, Cq7bx6, Zr7bx6, Zt7bx6, Zv7bx6, Zx7bx6, Zz7bx6, Z18bx6;
reg Z38bx6, Z58bx6, Z78bx6, Z98bx6, Zb8bx6, Zd8bx6, Zf8bx6, Zh8bx6, Zj8bx6, Zl8bx6;
reg Zn8bx6, Zp8bx6, Zr8bx6, Yt8bx6, Xv8bx6, Ux8bx6, Rz8bx6, N19bx6, J39bx6, F59bx6;
reg B79bx6, Q89bx6, Ua9bx6, Tc9bx6, Pe9bx6, Lg9bx6, Hi9bx6, Dk9bx6, Zl9bx6, Vn9bx6;
reg Jp9bx6, Lr9bx6, Nt9bx6, Nv9bx6, Ox9bx6, Pz9bx6, R1abx6, T3abx6, V5abx6, X7abx6;
reg Z9abx6, Bcabx6, Ceabx6, Ggabx6, Liabx6, Qkabx6, Nmabx6, Koabx6, Hqabx6, Esabx6;
reg Buabx6, Yvabx6, Nxabx6, Kzabx6, L1bbx6, L3bbx6, N5bbx6, P7bbx6, L9bbx6, Pbbbx6;
reg Pdbbx6, Ufbbx6, Lhbbx6, Qjbbx6, Nlbbx6, Knbbx6, Hpbbx6, Erbbx6, Btbbx6, Yubbx6;
reg Nwbbx6, Nybbx6, N0cbx6, S2cbx6, J4cbx6, A6cbx6, F8cbx6, Facbx6, Cccbx6, Zdcbx6;
reg Wfcbx6, Thcbx6, Qjcbx6, Nlcbx6, Cncbx6, Hpcbx6, Drcbx6, Itcbx6, Fvcbx6, Cxcbx6;
reg Zycbx6, W0dbx6, T2dbx6, Q4dbx6, F6dbx6, F8dbx6, Kadbx6, Bcdbx6, Sddbx6, Jfdbx6;
reg Ahdbx6, Fjdbx6, Fldbx6, Cndbx6, Zodbx6, Wqdbx6, Tsdbx6, Qudbx6, Nwdbx6, Cydbx6;
reg H0ebx6, M2ebx6, M4ebx6, J6ebx6, G8ebx6, Daebx6, Acebx6, Xdebx6, Ufebx6, Jhebx6;
reg Ojebx6, Tlebx6, Tnebx6, Tpebx6, Trebx6, Ttebx6, Tvebx6, Txebx6, Tzebx6, T1fbx6;
reg T3fbx6, T5fbx6, T7fbx6, T9fbx6, Tbfbx6, Tdfbx6, Tffbx6, Thfbx6, Tjfbx6, Qlfbx6;
reg Nnfbx6, Kpfbx6, Hrfbx6, Etfbx6, Bvfbx6, Qwfbx6, Vyfbx6, Y0gbx6, B3gbx6, C5gbx6;
reg D7gbx6, F9gbx6, Hbgbx6, Jdgbx6, Lfgbx6, Nhgbx6, Pjgbx6, Rlgbx6, Tngbx6, Vpgbx6;
reg Urgbx6, Ztgbx6, Zvgbx6, Wxgbx6, Tzgbx6, Q1hbx6, N3hbx6, K5hbx6, H7hbx6, W8hbx6;
reg Wahbx6, Tchbx6, Qehbx6, Eghbx6, Gihbx6, Ikhbx6, Imhbx6, Johbx6, Kqhbx6, Kshbx6;
reg Muhbx6, Owhbx6, Oyhbx6, P0ibx6, Q2ibx6, F4ibx6, X5ibx6, R7ibx6, R9ibx6, Rbibx6;
reg Rdibx6, Rfibx6, Rhibx6, Rjibx6, Rlibx6, Rnibx6, Rpibx6, Rribx6, Rtibx6, Rvibx6;
reg Qxibx6, Pzibx6, O1jbx6, N3jbx6, J5jbx6, F7jbx6, B9jbx6, Xajbx6, Tcjbx6, Pejbx6;
reg Pgjbx6, Rijbx6, Tkjbx6, Tmjbx6, Uojbx6, Vqjbx6, Usjbx6, Tujbx6, Swjbx6, Syjbx6;
reg S0kbx6, T2kbx6, S4kbx6, T6kbx6, T8kbx6, Qakbx6, Nckbx6, Rekbx6, Tgkbx6, Tikbx6;
reg Pkkbx6, Lmkbx6, Cokbx6, Dqkbx6;
wire [33:0] Vrkbx6;
wire [31:0] Ntkbx6;
wire [31:0] Nvkbx6;
wire [33:0] Nxkbx6;
wire [33:0] Ozkbx6;

assign HPROT[1] = 1'b1;
assign HBURST[2] = 1'b0;
assign HBURST[1] = 1'b0;
assign HBURST[0] = 1'b0;
assign HMASTLOCK = 1'b0;
assign HSIZE[2] = 1'b0;
assign HTRANS[0] = 1'b0;
assign nTDOEN = 1'b0;
assign WICENACK = 1'b0;
assign TDO = 1'b0;
assign WICSENSE[0] = 1'b0;
assign WICSENSE[1] = 1'b0;
assign WICSENSE[2] = 1'b0;
assign WICSENSE[3] = 1'b0;
assign WICSENSE[4] = 1'b0;
assign WICSENSE[5] = 1'b0;
assign WICSENSE[6] = 1'b0;
assign WICSENSE[7] = 1'b0;
assign WICSENSE[8] = 1'b0;
assign WICSENSE[9] = 1'b0;
assign WICSENSE[10] = 1'b0;
assign WICSENSE[11] = 1'b0;
assign WICSENSE[12] = 1'b0;
assign WICSENSE[13] = 1'b0;
assign WICSENSE[14] = 1'b0;
assign WICSENSE[15] = 1'b0;
assign WICSENSE[16] = 1'b0;
assign WICSENSE[17] = 1'b0;
assign WICSENSE[18] = 1'b0;
assign WICSENSE[19] = 1'b0;
assign WICSENSE[20] = 1'b0;
assign WICSENSE[21] = 1'b0;
assign WICSENSE[22] = 1'b0;
assign WICSENSE[23] = 1'b0;
assign WICSENSE[24] = 1'b0;
assign WICSENSE[25] = 1'b0;
assign WICSENSE[26] = 1'b0;
assign WICSENSE[27] = 1'b0;
assign WICSENSE[28] = 1'b0;
assign WICSENSE[29] = 1'b0;
assign WICSENSE[30] = 1'b0;
assign WICSENSE[31] = 1'b0;
assign WICSENSE[32] = 1'b0;
assign WICSENSE[33] = 1'b0;
assign WAKEUP = 1'b0;
assign Qmdhu6 = Evhpw6;
assign Pndhu6 = Hwhpw6;
assign Oodhu6 = Kxhpw6;
assign O5ohu6 = Nyhpw6;
assign Gwnhu6 = T0ipw6;
assign X0ohu6 = A3ipw6;
assign Q8nhu6 = A5ipw6;
assign Iahpw6[0] = W6ipw6;
assign Shhpw6[1] = M8ipw6;
assign Zvdpw6 = (!Qaipw6);
assign Odgpw6[30] = Tcipw6;
assign vis_r1_o[30] = Weipw6;
assign H8gpw6[0] = Wgipw6;
assign Ppfpw6[3] = Xiipw6;
assign D7fpw6[3] = Wkipw6;
assign X3fpw6[3] = Vmipw6;
assign vis_r11_o[30] = Uoipw6;
assign vis_r11_o[28] = Uqipw6;
assign Vbgpw6[28] = Usipw6;
assign vis_r11_o[4] = Vuipw6;
assign vis_r0_o[4] = Uwipw6;
assign Bagpw6[12] = Tyipw6;
assign Tzfpw6[12] = V0jpw6;
assign vis_r11_o[20] = X2jpw6;
assign vis_psp_o[18] = X4jpw6;
assign Bagpw6[20] = X6jpw6;
assign Tzfpw6[20] = Z8jpw6;
assign vis_r11_o[12] = Bbjpw6;
assign vis_psp_o[10] = Bdjpw6;
assign vis_apsr_o[2] = Bfjpw6;
assign H6ghu6 = Vgjpw6;
assign vis_apsr_o[1] = Qijpw6;
assign vis_r11_o[29] = Kkjpw6;
assign vis_r8_o[29] = Kmjpw6;
assign Vbgpw6[29] = Kojpw6;
assign vis_pc_o[28] = Lqjpw6;
assign Vchhu6 = Isjpw6;
assign Cyfpw6[6] = Aujpw6;
assign Cyfpw6[7] = Yvjpw6;
assign H2fpw6[1] = Wxjpw6;
assign Ivfhu6 = Vzjpw6;
assign S8fpw6[3] = U1kpw6;
assign vis_r11_o[5] = T3kpw6;
assign vis_r8_o[5] = S5kpw6;
assign Bagpw6[13] = R7kpw6;
assign Tzfpw6[13] = T9kpw6;
assign vis_ipsr_o[5] = Vbkpw6;
assign vis_r11_o[21] = Rdkpw6;
assign vis_psp_o[19] = Rfkpw6;
assign Bagpw6[21] = Rhkpw6;
assign Tzfpw6[21] = Tjkpw6;
assign vis_r11_o[13] = Vlkpw6;
assign vis_psp_o[11] = Vnkpw6;
assign Hwmhu6 = Vpkpw6;
assign Uthpw6[24] = Nrkpw6;
assign Iahpw6[23] = Stkpw6;
assign Shhpw6[24] = Jvkpw6;
assign Vbgpw6[24] = Oxkpw6;
assign vis_tbit_o = Pzkpw6;
assign Fkfpw6[0] = I1lpw6;
assign Uthpw6[0] = H3lpw6;
assign Tonhu6 = L5lpw6;
assign Yenhu6 = B7lpw6;
assign Hknhu6 = Y8lpw6;
assign Ighpw6[2] = Kalpw6;
assign Ighpw6[0] = Bclpw6;
assign Ighpw6[1] = Sdlpw6;
assign Ighpw6[3] = Jflpw6;
assign Fnnhu6 = Ahlpw6;
assign Mdhpw6[3] = Rilpw6;
assign Ighpw6[4] = Yklpw6;
assign Ighpw6[5] = Pmlpw6;
assign Mdhpw6[2] = Golpw6;
assign Mdhpw6[1] = Vplpw6;
assign Mdhpw6[0] = Krlpw6;
assign Ulnhu6 = Zslpw6;
assign Pinhu6 = Oulpw6;
assign B7nhu6 = Kwlpw6;
assign Ubnhu6 = Gylpw6;
assign Iahpw6[6] = Yzlpw6;
assign Shhpw6[7] = O1mpw6;
assign R4gpw6[9] = S3mpw6;
assign Ppfpw6[1] = T5mpw6;
assign D7fpw6[1] = S7mpw6;
assign S8fpw6[1] = R9mpw6;
assign vis_r11_o[3] = Qbmpw6;
assign vis_r8_o[3] = Pdmpw6;
assign Bagpw6[11] = Ofmpw6;
assign vis_ipsr_o[3] = Qhmpw6;
assign vis_r11_o[27] = Mjmpw6;
assign vis_r8_o[27] = Mlmpw6;
assign Ikghu6 = Mnmpw6;
assign Ppfpw6[2] = Jpmpw6;
assign D7fpw6[2] = Irmpw6;
assign X3fpw6[2] = Htmpw6;
assign vis_r0_o[30] = Gvmpw6;
assign vis_r0_o[3] = Gxmpw6;
assign vis_r0_o[5] = Fzmpw6;
assign vis_r0_o[27] = E1npw6;
assign vis_r0_o[29] = E3npw6;
assign vis_r0_o[21] = E5npw6;
assign vis_r0_o[20] = E7npw6;
assign vis_r0_o[13] = E9npw6;
assign vis_r0_o[12] = Ebnpw6;
assign vis_r0_o[28] = Ednpw6;
assign vis_r11_o[31] = Efnpw6;
assign vis_r0_o[31] = Ehnpw6;
assign vis_r1_o[31] = Ejnpw6;
assign H8gpw6[1] = Elnpw6;
assign Stdhu6 = Fnnpw6;
assign E5ehu6 = Fpnpw6;
assign vis_apsr_o[3] = Arnpw6;
assign Fkfpw6[31] = Usnpw6;
assign Uthpw6[31] = Uunpw6;
assign Iahpw6[30] = Zwnpw6;
assign Vmdpw6 = (!Qynpw6);
assign Fanhu6 = I0opw6;
assign Iahpw6[4] = D2opw6;
assign Shhpw6[5] = T3opw6;
assign Bagpw6[5] = X5opw6;
assign Tzfpw6[5] = Y7opw6;
assign Fsdhu6 = Z9opw6;
assign SLEEPHOLDACKn = Xbopw6;
assign E6phu6 = (!Xbopw6);
assign C0ehu6 = Ydopw6;
assign Cyfpw6[3] = Ufopw6;
assign H2fpw6[0] = Shopw6;
assign vis_r9_o[4] = Rjopw6;
assign vis_r9_o[30] = Qlopw6;
assign vis_r9_o[31] = Qnopw6;
assign vis_r9_o[3] = Qpopw6;
assign vis_r9_o[5] = Propw6;
assign vis_r9_o[27] = Otopw6;
assign vis_r9_o[29] = Ovopw6;
assign vis_r9_o[21] = Oxopw6;
assign vis_r9_o[20] = Ozopw6;
assign vis_r9_o[13] = O1ppw6;
assign vis_r9_o[12] = O3ppw6;
assign vis_r5_o[4] = O5ppw6;
assign vis_r5_o[30] = N7ppw6;
assign vis_r5_o[31] = N9ppw6;
assign vis_r5_o[3] = Nbppw6;
assign vis_r5_o[5] = Mdppw6;
assign vis_r5_o[27] = Lfppw6;
assign vis_r5_o[29] = Lhppw6;
assign vis_r5_o[21] = Ljppw6;
assign vis_r5_o[20] = Llppw6;
assign vis_r5_o[13] = Lnppw6;
assign vis_r5_o[12] = Lpppw6;
assign vis_r1_o[4] = Lrppw6;
assign vis_r1_o[3] = Ktppw6;
assign vis_r1_o[5] = Jvppw6;
assign vis_r1_o[27] = Ixppw6;
assign vis_r1_o[29] = Izppw6;
assign vis_r1_o[21] = I1qpw6;
assign vis_r1_o[20] = I3qpw6;
assign vis_r1_o[13] = I5qpw6;
assign vis_r1_o[12] = I7qpw6;
assign vis_r1_o[28] = I9qpw6;
assign Fkfpw6[28] = Ibqpw6;
assign Uthpw6[28] = Idqpw6;
assign Iahpw6[27] = Nfqpw6;
assign Zbhpw6[28] = Ehqpw6;
assign Punhu6 = Cjqpw6;
assign CDBGPWRUPREQ = Xkqpw6;
assign W9ohu6 = (!Xkqpw6);
assign Iqnhu6 = Gnqpw6;
assign Cjhpw6[0] = Gpqpw6;
assign Cjhpw6[1] = Nrqpw6;
assign G2ohu6 = Utqpw6;
assign Q7ohu6 = Xvqpw6;
assign Lznhu6 = Xxqpw6;
assign Shhpw6[31] = Yzqpw6;
assign Shhpw6[28] = D2rpw6;
assign Shhpw6[0] = I4rpw6;
assign Bagpw6[0] = M6rpw6;
assign Tzfpw6[0] = N8rpw6;
assign Tzfpw6[1] = Oarpw6;
assign vis_ipsr_o[1] = Pcrpw6;
assign vis_pc_o[0] = Lerpw6;
assign S1ehu6 = Hgrpw6;
assign H4ghu6 = Hirpw6;
assign S8fpw6[5] = Fkrpw6;
assign vis_r0_o[7] = Emrpw6;
assign vis_r1_o[7] = Dorpw6;
assign vis_r9_o[7] = Cqrpw6;
assign vis_r11_o[7] = Bsrpw6;
assign vis_r5_o[7] = Aurpw6;
assign vis_r8_o[7] = Zvrpw6;
assign Odgpw6[15] = Yxrpw6;
assign vis_r0_o[6] = B0spw6;
assign vis_r1_o[6] = A2spw6;
assign vis_r9_o[6] = Z3spw6;
assign vis_r11_o[6] = Y5spw6;
assign vis_r5_o[6] = X7spw6;
assign vis_r8_o[6] = W9spw6;
assign R4gpw6[10] = Vbspw6;
assign Ppfpw6[0] = Xdspw6;
assign D7fpw6[0] = Wfspw6;
assign X3fpw6[0] = Vhspw6;
assign Bagpw6[16] = Ujspw6;
assign Tzfpw6[16] = Wlspw6;
assign vis_r0_o[24] = Ynspw6;
assign vis_r1_o[24] = Ypspw6;
assign vis_r9_o[24] = Yrspw6;
assign vis_r11_o[24] = Ytspw6;
assign vis_r5_o[24] = Yvspw6;
assign vis_r8_o[24] = Yxspw6;
assign Jfgpw6[0] = Yzspw6;
assign vis_r0_o[25] = Z1tpw6;
assign vis_r1_o[25] = Z3tpw6;
assign vis_r9_o[25] = Z5tpw6;
assign vis_r11_o[25] = Z7tpw6;
assign vis_r5_o[25] = Z9tpw6;
assign vis_psp_o[23] = Zbtpw6;
assign Yyghu6 = Zdtpw6;
assign vis_r9_o[2] = Yftpw6;
assign vis_r11_o[2] = Xhtpw6;
assign vis_r5_o[2] = Wjtpw6;
assign vis_r0_o[2] = Vltpw6;
assign vis_r1_o[2] = Untpw6;
assign Bagpw6[10] = Tptpw6;
assign Tzfpw6[10] = Vrtpw6;
assign vis_r0_o[26] = Xttpw6;
assign vis_r1_o[26] = Xvtpw6;
assign vis_r9_o[26] = Xxtpw6;
assign vis_r11_o[26] = Xztpw6;
assign vis_r5_o[26] = X1upw6;
assign vis_r8_o[26] = X3upw6;
assign Vbgpw6[26] = X5upw6;
assign vis_r0_o[17] = Y7upw6;
assign vis_r1_o[17] = Y9upw6;
assign vis_r9_o[17] = Ybupw6;
assign vis_r11_o[17] = Ydupw6;
assign vis_r5_o[17] = Yfupw6;
assign vis_psp_o[15] = Yhupw6;
assign Bagpw6[17] = Yjupw6;
assign Tzfpw6[17] = Amupw6;
assign Tzfpw6[23] = Coupw6;
assign vis_pc_o[6] = Equpw6;
assign Fkfpw6[7] = Asupw6;
assign Jfgpw6[4] = Ztupw6;
assign vis_pc_o[30] = Awupw6;
assign Cyfpw6[1] = Xxupw6;
assign Cyfpw6[0] = Vzupw6;
assign Cyfpw6[4] = T1vpw6;
assign Cyfpw6[5] = R3vpw6;
assign Y7ghu6 = P5vpw6;
assign DBGRESTARTED = K7vpw6;
assign Daohu6 = (!K7vpw6);
assign V9ghu6 = F9vpw6;
assign Uthpw6[19] = Gbvpw6;
assign Iahpw6[18] = Ldvpw6;
assign Shhpw6[19] = Cfvpw6;
assign Bagpw6[19] = Hhvpw6;
assign vis_r0_o[19] = Jjvpw6;
assign vis_r1_o[19] = Jlvpw6;
assign vis_r9_o[19] = Jnvpw6;
assign vis_r11_o[19] = Jpvpw6;
assign vis_r5_o[19] = Jrvpw6;
assign vis_psp_o[17] = Jtvpw6;
assign Svdpw6 = (!Jvvpw6);
assign D7fpw6[14] = Dxvpw6;
assign H2fpw6[2] = Dzvpw6;
assign Npdhu6 = C1wpw6;
assign Vbgpw6[0] = C3wpw6;
assign vis_r0_o[16] = C5wpw6;
assign vis_r1_o[16] = C7wpw6;
assign vis_r9_o[16] = C9wpw6;
assign vis_r11_o[16] = Cbwpw6;
assign vis_r5_o[16] = Cdwpw6;
assign vis_psp_o[14] = Cfwpw6;
assign Fkfpw6[16] = Chwpw6;
assign Uthpw6[16] = Cjwpw6;
assign Iahpw6[15] = Hlwpw6;
assign Shhpw6[16] = Ymwpw6;
assign Jshpw6[16] = Dpwpw6;
assign X8hpw6[6] = Sqwpw6;
assign Uthpw6[18] = Kswpw6;
assign Iahpw6[17] = Puwpw6;
assign Shhpw6[18] = Gwwpw6;
assign Bagpw6[18] = Lywpw6;
assign Tzfpw6[18] = N0xpw6;
assign vis_r0_o[18] = P2xpw6;
assign vis_r1_o[18] = P4xpw6;
assign vis_r9_o[18] = P6xpw6;
assign vis_r11_o[18] = P8xpw6;
assign vis_r5_o[18] = Paxpw6;
assign vis_psp_o[16] = Pcxpw6;
assign Aghhu6 = Pexpw6;
assign D7fpw6[4] = Jgxpw6;
assign X3fpw6[1] = Iixpw6;
assign vis_r0_o[10] = Hkxpw6;
assign vis_r1_o[10] = Hmxpw6;
assign vis_r9_o[10] = Hoxpw6;
assign vis_r11_o[10] = Hqxpw6;
assign vis_r5_o[10] = Hsxpw6;
assign vis_psp_o[8] = Huxpw6;
assign Fkfpw6[10] = Gwxpw6;
assign Uthpw6[10] = Gyxpw6;
assign Iahpw6[9] = L0ypw6;
assign Shhpw6[10] = C2ypw6;
assign Jshpw6[10] = H4ypw6;
assign Jfgpw6[2] = W5ypw6;
assign Ntfhu6 = X7ypw6;
assign D7fpw6[15] = U9ypw6;
assign S8fpw6[4] = Ubypw6;
assign vis_r0_o[1] = Tdypw6;
assign vis_r1_o[1] = Sfypw6;
assign vis_r9_o[1] = Rhypw6;
assign vis_r11_o[1] = Qjypw6;
assign vis_r5_o[1] = Plypw6;
assign vis_r14_o[1] = Onypw6;
assign vis_control_o = Npypw6;
assign Vrfhu6 = Jrypw6;
assign vis_psp_o[0] = Ftypw6;
assign vis_psp_o[29] = Evypw6;
assign vis_psp_o[28] = Exypw6;
assign vis_psp_o[2] = Ezypw6;
assign vis_psp_o[1] = D1zpw6;
assign vis_psp_o[3] = C3zpw6;
assign vis_psp_o[4] = B5zpw6;
assign vis_psp_o[5] = A7zpw6;
assign vis_psp_o[22] = Z8zpw6;
assign vis_psp_o[24] = Zazpw6;
assign vis_psp_o[25] = Zczpw6;
assign vis_psp_o[27] = Zezpw6;
assign vis_msp_o[0] = Zgzpw6;
assign vis_msp_o[29] = Yizpw6;
assign vis_msp_o[28] = Ykzpw6;
assign vis_msp_o[2] = Ymzpw6;
assign vis_msp_o[1] = Xozpw6;
assign vis_msp_o[3] = Wqzpw6;
assign vis_msp_o[4] = Vszpw6;
assign vis_msp_o[5] = Uuzpw6;
assign vis_msp_o[22] = Twzpw6;
assign vis_msp_o[24] = Tyzpw6;
assign vis_msp_o[25] = T00qw6;
assign vis_msp_o[27] = T20qw6;
assign vis_msp_o[23] = T40qw6;
assign vis_msp_o[19] = T60qw6;
assign vis_msp_o[18] = T80qw6;
assign vis_msp_o[17] = Ta0qw6;
assign vis_msp_o[16] = Tc0qw6;
assign vis_msp_o[15] = Te0qw6;
assign vis_msp_o[14] = Tg0qw6;
assign vis_msp_o[11] = Ti0qw6;
assign vis_msp_o[10] = Tk0qw6;
assign vis_msp_o[8] = Tm0qw6;
assign vis_msp_o[6] = So0qw6;
assign Bagpw6[8] = Rq0qw6;
assign Tzfpw6[8] = Ss0qw6;
assign vis_r0_o[8] = Tu0qw6;
assign vis_r1_o[8] = Sw0qw6;
assign vis_r9_o[8] = Ry0qw6;
assign vis_r11_o[8] = Q01qw6;
assign vis_r5_o[8] = P21qw6;
assign vis_psp_o[6] = O41qw6;
assign Fkfpw6[8] = N61qw6;
assign Uthpw6[8] = M81qw6;
assign Iahpw6[7] = Qa1qw6;
assign Shhpw6[8] = Gc1qw6;
assign Jshpw6[8] = Ke1qw6;
assign Jshpw6[9] = Yf1qw6;
assign Uthpw6[9] = Mh1qw6;
assign Iahpw6[8] = Qj1qw6;
assign Shhpw6[9] = Gl1qw6;
assign Fkfpw6[9] = Kn1qw6;
assign vis_r0_o[9] = Jp1qw6;
assign vis_r1_o[9] = Ir1qw6;
assign vis_r9_o[9] = Ht1qw6;
assign vis_r11_o[9] = Gv1qw6;
assign vis_r5_o[9] = Fx1qw6;
assign vis_r7_o[9] = Ez1qw6;
assign vis_pc_o[27] = D12qw6;
assign vis_pc_o[29] = A32qw6;
assign Uthpw6[30] = X42qw6;
assign Iahpw6[29] = C72qw6;
assign Zbhpw6[30] = T82qw6;
assign Shhpw6[30] = Ra2qw6;
assign Jshpw6[30] = Wc2qw6;
assign X8hpw6[1] = Le2qw6;
assign A2nhu6 = Dg2qw6;
assign R6hhu6 = Uh2qw6;
assign D8hhu6 = Nj2qw6;
assign Uthpw6[25] = Fl2qw6;
assign Iahpw6[24] = Kn2qw6;
assign Shhpw6[25] = Bp2qw6;
assign Jehhu6 = Gr2qw6;
assign P9hhu6 = Bt2qw6;
assign Uthpw6[3] = Xu2qw6;
assign Iahpw6[2] = Bx2qw6;
assign Jdnhu6 = Ry2qw6;
assign Shhpw6[3] = L03qw6;
assign Tnhpw6[3] = P23qw6;
assign X8hpw6[3] = D43qw6;
assign Uthpw6[4] = V53qw6;
assign Iahpw6[3] = Z73qw6;
assign Shhpw6[4] = P93qw6;
assign Cynhu6 = Tb3qw6;
assign Jshpw6[7] = Nd3qw6;
assign Jshpw6[5] = Bf3qw6;
assign Jshpw6[4] = Pg3qw6;
assign X8hpw6[4] = Di3qw6;
assign Tnhpw6[1] = Vj3qw6;
assign Jshpw6[18] = Jl3qw6;
assign Jshpw6[19] = Ym3qw6;
assign Jshpw6[24] = No3qw6;
assign Jshpw6[29] = Cq3qw6;
assign Uthpw6[29] = Rr3qw6;
assign Iahpw6[28] = Wt3qw6;
assign Shhpw6[29] = Nv3qw6;
assign Fkfpw6[29] = Sx3qw6;
assign Yyfhu6 = Sz3qw6;
assign D7fpw6[13] = P14qw6;
assign vis_r9_o[23] = P34qw6;
assign vis_r11_o[23] = P54qw6;
assign vis_msp_o[21] = Gp6ax6;
assign vis_psp_o[21] = Gr6ax6;
assign vis_r5_o[23] = Gt6ax6;
assign vis_r0_o[23] = Gv6ax6;
assign vis_r1_o[23] = Gx6ax6;
assign L1gpw6[1] = Gz6ax6;
assign Zlghu6 = F17ax6;
assign vis_pc_o[22] = C37ax6;
assign Fkfpw6[15] = Z47ax6;
assign Uthpw6[15] = Z67ax6;
assign Iahpw6[14] = E97ax6;
assign Shhpw6[15] = Va7ax6;
assign Jshpw6[15] = Ad7ax6;
assign X8hpw6[2] = Pe7ax6;
assign Uthpw6[2] = Hg7ax6;
assign Iahpw6[1] = Li7ax6;
assign Shhpw6[2] = Bk7ax6;
assign Hbhhu6 = Fm7ax6;
assign Tnhpw6[2] = Xn7ax6;
assign Ftghu6 = Lp7ax6;
assign Tzfpw6[19] = Nr7ax6;
assign Tzfpw6[11] = Pt7ax6;
assign Tzfpw6[6] = Rv7ax6;
assign vis_r0_o[14] = Sx7ax6;
assign vis_r1_o[14] = Sz7ax6;
assign vis_r9_o[14] = S18ax6;
assign vis_r11_o[14] = S38ax6;
assign vis_r5_o[14] = S58ax6;
assign vis_msp_o[12] = S78ax6;
assign vis_psp_o[12] = S98ax6;
assign Fkfpw6[14] = Sb8ax6;
assign Uthpw6[14] = Sd8ax6;
assign Iahpw6[13] = Xf8ax6;
assign Iahpw6[12] = Oh8ax6;
assign Shhpw6[13] = Fj8ax6;
assign Jshpw6[13] = Kl8ax6;
assign X8hpw6[5] = Zm8ax6;
assign Uthpw6[12] = Ro8ax6;
assign Iahpw6[11] = Wq8ax6;
assign Shhpw6[12] = Ns8ax6;
assign Jshpw6[12] = Su8ax6;
assign X8hpw6[0] = Hw8ax6;
assign Lwgpw6[0] = Zx8ax6;
assign Lwgpw6[2] = Vz8ax6;
assign Lwgpw6[1] = R19ax6;
assign V5hpw6[0] = N39ax6;
assign K7hpw6[30] = J59ax6;
assign K7hpw6[25] = G79ax6;
assign K7hpw6[24] = D99ax6;
assign K7hpw6[19] = Ab9ax6;
assign K7hpw6[18] = Xc9ax6;
assign K7hpw6[16] = Ue9ax6;
assign K7hpw6[15] = Rg9ax6;
assign K7hpw6[13] = Oi9ax6;
assign K7hpw6[12] = Lk9ax6;
assign K7hpw6[10] = Im9ax6;
assign K7hpw6[8] = Fo9ax6;
assign K7hpw6[7] = Bq9ax6;
assign K7hpw6[5] = Xr9ax6;
assign K7hpw6[4] = Tt9ax6;
assign K7hpw6[3] = Pv9ax6;
assign K7hpw6[2] = Lx9ax6;
assign V5hpw6[1] = Hz9ax6;
assign Pzgpw6[0] = D1aax6;
assign E1hpw6[30] = Z2aax6;
assign E1hpw6[25] = W4aax6;
assign E1hpw6[24] = T6aax6;
assign E1hpw6[19] = Q8aax6;
assign E1hpw6[18] = Naaax6;
assign E1hpw6[16] = Kcaax6;
assign E1hpw6[15] = Heaax6;
assign E1hpw6[13] = Egaax6;
assign E1hpw6[12] = Biaax6;
assign E1hpw6[10] = Yjaax6;
assign E1hpw6[8] = Vlaax6;
assign E1hpw6[7] = Rnaax6;
assign E1hpw6[5] = Npaax6;
assign E1hpw6[4] = Jraax6;
assign E1hpw6[3] = Ftaax6;
assign E1hpw6[2] = Bvaax6;
assign Pzgpw6[1] = Xwaax6;
assign R2hpw6[0] = Tyaax6;
assign R2hpw6[2] = P0bax6;
assign R2hpw6[1] = L2bax6;
assign Kohhu6 = H4bax6;
assign G4hpw6[1] = X5bax6;
assign G4hpw6[2] = T7bax6;
assign G4hpw6[3] = P9bax6;
assign G4hpw6[4] = Lbbax6;
assign Aygpw6[1] = Hdbax6;
assign Aygpw6[2] = Dfbax6;
assign Aygpw6[3] = Zgbax6;
assign Aygpw6[4] = Vibax6;
assign Dhgpw6[2] = Rkbax6;
assign Dhgpw6[4] = Hmbax6;
assign Dhgpw6[1] = Xnbax6;
assign Gtgpw6[2] = Opbax6;
assign Engpw6[27] = Krbax6;
assign Gtgpw6[25] = Htbax6;
assign Gtgpw6[24] = Evbax6;
assign Gtgpw6[19] = Bxbax6;
assign Gtgpw6[18] = Yybax6;
assign Gtgpw6[16] = V0cax6;
assign Gtgpw6[15] = S2cax6;
assign Gtgpw6[13] = P4cax6;
assign Gtgpw6[12] = M6cax6;
assign Gtgpw6[10] = J8cax6;
assign Gtgpw6[8] = Facax6;
assign Gtgpw6[7] = Bccax6;
assign Gtgpw6[5] = Xdcax6;
assign Gtgpw6[4] = Tfcax6;
assign Gtgpw6[3] = Phcax6;
assign Smhhu6 = Ljcax6;
assign Togpw6[2] = Hlcax6;
assign Ligpw6[27] = Dncax6;
assign Togpw6[25] = Apcax6;
assign Togpw6[24] = Xqcax6;
assign Togpw6[19] = Uscax6;
assign Togpw6[18] = Rucax6;
assign Togpw6[16] = Owcax6;
assign Togpw6[15] = Lycax6;
assign Togpw6[13] = I0dax6;
assign Togpw6[12] = F2dax6;
assign Togpw6[10] = C4dax6;
assign Togpw6[8] = Y5dax6;
assign Togpw6[7] = U7dax6;
assign Togpw6[5] = Q9dax6;
assign Togpw6[4] = Mbdax6;
assign Togpw6[3] = Iddax6;
assign Qhhhu6 = Efdax6;
assign Gqgpw6[2] = Ahdax6;
assign Akgpw6[27] = Widax6;
assign Gqgpw6[25] = Tkdax6;
assign Gqgpw6[24] = Qmdax6;
assign Gqgpw6[19] = Nodax6;
assign Gqgpw6[18] = Kqdax6;
assign Gqgpw6[16] = Hsdax6;
assign Gqgpw6[15] = Eudax6;
assign Gqgpw6[13] = Bwdax6;
assign Gqgpw6[12] = Yxdax6;
assign Gqgpw6[10] = Vzdax6;
assign Gqgpw6[8] = R1eax6;
assign Gqgpw6[7] = N3eax6;
assign Gqgpw6[5] = J5eax6;
assign Gqgpw6[4] = F7eax6;
assign Gqgpw6[3] = B9eax6;
assign Ijhhu6 = Xaeax6;
assign Trgpw6[2] = Tceax6;
assign Plgpw6[27] = Peeax6;
assign Trgpw6[25] = Mgeax6;
assign Trgpw6[24] = Jieax6;
assign Trgpw6[19] = Gkeax6;
assign Trgpw6[18] = Dmeax6;
assign Trgpw6[16] = Aoeax6;
assign Trgpw6[15] = Xpeax6;
assign Trgpw6[13] = Ureax6;
assign Trgpw6[12] = Rteax6;
assign Trgpw6[10] = Oveax6;
assign Trgpw6[8] = Kxeax6;
assign Trgpw6[7] = Gzeax6;
assign Trgpw6[5] = C1fax6;
assign Trgpw6[4] = Y2fax6;
assign Trgpw6[3] = U4fax6;
assign Alhhu6 = Q6fax6;
assign T0hhu6 = M8fax6;
assign H2hhu6 = Eafax6;
assign E5hhu6 = Sbfax6;
assign S3hhu6 = Hdfax6;
assign Uthpw6[6] = Vefax6;
assign Iahpw6[5] = Zgfax6;
assign Omdpw6 = (!Pifax6);
assign N3nhu6 = Okfax6;
assign Cjhpw6[2] = Nmfax6;
assign Sqhpw6[1] = Uofax6;
assign Sqhpw6[0] = Sqfax6;
assign Dtnhu6 = Qsfax6;
assign S3ohu6 = Qufax6;
assign Rrnhu6 = Qwfax6;
assign Rgnhu6 = Ryfax6;
assign Cjhpw6[3] = J0gax6;
assign K7hpw6[31] = Q2gax6;
assign E1hpw6[31] = N4gax6;
assign Engpw6[28] = K6gax6;
assign Plgpw6[28] = H8gax6;
assign Akgpw6[28] = Eagax6;
assign Ligpw6[28] = Bcgax6;
assign Jshpw6[31] = Ydgax6;
assign K7hpw6[28] = Nfgax6;
assign E1hpw6[28] = Khgax6;
assign Gtgpw6[28] = Hjgax6;
assign Trgpw6[28] = Elgax6;
assign Gqgpw6[28] = Bngax6;
assign Togpw6[28] = Yogax6;
assign Jshpw6[28] = Vqgax6;
assign Aphpw6[1] = Ksgax6;
assign Aphpw6[2] = Dugax6;
assign R0nhu6 = Wvgax6;
assign Jzmhu6 = Jxgax6;
assign Sbghu6 = Vygax6;
assign vis_pc_o[26] = U0hax6;
assign vis_pc_o[25] = R2hax6;
assign vis_pc_o[24] = O4hax6;
assign vis_pc_o[23] = L6hax6;
assign vis_pc_o[20] = I8hax6;
assign vis_pc_o[19] = Fahax6;
assign vis_pc_o[18] = Cchax6;
assign vis_pc_o[17] = Zdhax6;
assign vis_pc_o[16] = Wfhax6;
assign vis_pc_o[15] = Thhax6;
assign vis_pc_o[13] = Qjhax6;
assign vis_pc_o[12] = Nlhax6;
assign vis_pc_o[11] = Knhax6;
assign vis_pc_o[7] = Hphax6;
assign vis_pc_o[5] = Drhax6;
assign vis_pc_o[4] = Zshax6;
assign vis_pc_o[3] = Vuhax6;
assign vis_pc_o[2] = Rwhax6;
assign vis_pc_o[1] = Nyhax6;
assign Sufpw6[1] = J0iax6;
assign Ppfpw6[4] = G2iax6;
assign Ppfpw6[5] = F4iax6;
assign Ppfpw6[14] = E6iax6;
assign Ppfpw6[6] = E8iax6;
assign N2ghu6 = Daiax6;
assign Fvdhu6 = Bciax6;
assign T6ehu6 = Zdiax6;
assign vis_primask_o = Xfiax6;
assign Dhgpw6[3] = Thiax6;
assign vis_ipsr_o[4] = Ijiax6;
assign vis_ipsr_o[0] = Eliax6;
assign vis_ipsr_o[2] = Aniax6;
assign Lvdpw6 = (!Woiax6);
assign Ppfpw6[7] = Zqiax6;
assign Ppfpw6[8] = Ysiax6;
assign Ppfpw6[9] = Xuiax6;
assign Ppfpw6[10] = Wwiax6;
assign Ppfpw6[11] = Wyiax6;
assign Ppfpw6[12] = W0jax6;
assign Ppfpw6[13] = W2jax6;
assign D7fpw6[6] = W4jax6;
assign S8fpw6[7] = V6jax6;
assign Dxfhu6 = U8jax6;
assign Hrfpw6[16] = Tajax6;
assign Hrfpw6[0] = Tcjax6;
assign Hrfpw6[15] = Sejax6;
assign Hrfpw6[13] = Sgjax6;
assign Hrfpw6[12] = Sijax6;
assign D7fpw6[12] = Skjax6;
assign Hrfpw6[11] = Smjax6;
assign D7fpw6[11] = Sojax6;
assign Hrfpw6[10] = Sqjax6;
assign D7fpw6[10] = Ssjax6;
assign Hrfpw6[9] = Sujax6;
assign D7fpw6[9] = Rwjax6;
assign Hrfpw6[8] = Qyjax6;
assign D7fpw6[8] = P0kax6;
assign Hrfpw6[7] = O2kax6;
assign D7fpw6[7] = N4kax6;
assign H2fpw6[3] = M6kax6;
assign Hrfpw6[6] = L8kax6;
assign Hrfpw6[5] = Kakax6;
assign D7fpw6[5] = Jckax6;
assign S8fpw6[8] = Iekax6;
assign S8fpw6[9] = Lgkax6;
assign S8fpw6[10] = Oikax6;
assign S8fpw6[11] = Rkkax6;
assign S8fpw6[6] = Umkax6;
assign Hrfpw6[4] = Tokax6;
assign S8fpw6[0] = Sqkax6;
assign S8fpw6[2] = Rskax6;
assign vis_r9_o[0] = Qukax6;
assign vis_r11_o[0] = Pwkax6;
assign vis_r5_o[0] = Oykax6;
assign vis_r0_o[0] = N0lax6;
assign vis_r1_o[0] = M2lax6;
assign Ppfpw6[16] = L4lax6;
assign Sufpw6[0] = L6lax6;
assign L3ehu6 = I8lax6;
assign Qwdhu6 = Halax6;
assign vis_r10_o[2] = Eclax6;
assign vis_r10_o[4] = Delax6;
assign vis_r10_o[23] = Cglax6;
assign vis_r10_o[30] = Cilax6;
assign vis_r10_o[31] = Cklax6;
assign vis_r10_o[0] = Cmlax6;
assign vis_r10_o[3] = Bolax6;
assign vis_r10_o[5] = Aqlax6;
assign vis_r10_o[6] = Zrlax6;
assign vis_r10_o[7] = Ytlax6;
assign vis_r10_o[24] = Xvlax6;
assign vis_r10_o[26] = Xxlax6;
assign vis_r10_o[27] = Xzlax6;
assign vis_r10_o[29] = X1max6;
assign vis_r10_o[1] = X3max6;
assign vis_r10_o[25] = W5max6;
assign vis_r10_o[21] = W7max6;
assign vis_r10_o[20] = W9max6;
assign vis_r10_o[19] = Wbmax6;
assign vis_r10_o[18] = Wdmax6;
assign vis_r10_o[17] = Wfmax6;
assign vis_r10_o[16] = Whmax6;
assign vis_r10_o[14] = Wjmax6;
assign vis_r10_o[13] = Wlmax6;
assign vis_r10_o[12] = Wnmax6;
assign vis_r10_o[10] = Wpmax6;
assign vis_r10_o[9] = Wrmax6;
assign vis_r10_o[8] = Vtmax6;
assign vis_r14_o[2] = Uvmax6;
assign vis_r14_o[4] = Txmax6;
assign vis_r14_o[23] = Szmax6;
assign vis_r14_o[30] = S1nax6;
assign vis_r14_o[31] = S3nax6;
assign vis_r14_o[0] = S5nax6;
assign vis_r14_o[3] = R7nax6;
assign vis_r14_o[5] = Q9nax6;
assign vis_r14_o[6] = Pbnax6;
assign vis_r14_o[7] = Odnax6;
assign vis_r14_o[24] = Nfnax6;
assign vis_r14_o[26] = Nhnax6;
assign vis_r14_o[27] = Njnax6;
assign vis_r14_o[29] = Nlnax6;
assign vis_r14_o[25] = Nnnax6;
assign vis_r14_o[21] = Npnax6;
assign vis_r14_o[20] = Nrnax6;
assign vis_r14_o[19] = Ntnax6;
assign vis_r14_o[18] = Nvnax6;
assign vis_r14_o[17] = Nxnax6;
assign vis_r14_o[16] = Nznax6;
assign vis_r14_o[14] = N1oax6;
assign vis_r14_o[13] = N3oax6;
assign vis_r14_o[12] = N5oax6;
assign vis_r14_o[10] = N7oax6;
assign vis_r14_o[8] = N9oax6;
assign vis_r6_o[2] = Mboax6;
assign vis_r6_o[4] = Ldoax6;
assign vis_r6_o[23] = Kfoax6;
assign vis_r6_o[30] = Khoax6;
assign vis_r6_o[31] = Kjoax6;
assign vis_r6_o[0] = Kloax6;
assign vis_r6_o[3] = Jnoax6;
assign vis_r6_o[5] = Ipoax6;
assign vis_r6_o[6] = Hroax6;
assign vis_r6_o[7] = Gtoax6;
assign vis_r6_o[24] = Fvoax6;
assign vis_r6_o[26] = Fxoax6;
assign vis_r6_o[27] = Fzoax6;
assign vis_r6_o[29] = F1pax6;
assign vis_r6_o[1] = F3pax6;
assign vis_r6_o[25] = E5pax6;
assign vis_r6_o[21] = E7pax6;
assign vis_r6_o[20] = E9pax6;
assign vis_r6_o[19] = Ebpax6;
assign vis_r6_o[18] = Edpax6;
assign vis_r6_o[17] = Efpax6;
assign vis_r6_o[16] = Ehpax6;
assign vis_r6_o[14] = Ejpax6;
assign vis_r6_o[13] = Elpax6;
assign vis_r6_o[12] = Enpax6;
assign vis_r6_o[10] = Eppax6;
assign vis_r6_o[9] = Erpax6;
assign vis_r6_o[8] = Dtpax6;
assign vis_r2_o[2] = Cvpax6;
assign vis_r2_o[4] = Bxpax6;
assign vis_r2_o[23] = Azpax6;
assign vis_r2_o[30] = A1qax6;
assign vis_r2_o[31] = A3qax6;
assign vis_r2_o[0] = A5qax6;
assign vis_r2_o[3] = Z6qax6;
assign vis_r2_o[5] = Y8qax6;
assign vis_r2_o[6] = Xaqax6;
assign vis_r2_o[7] = Wcqax6;
assign vis_r2_o[24] = Veqax6;
assign vis_r2_o[26] = Vgqax6;
assign vis_r2_o[27] = Viqax6;
assign vis_r2_o[29] = Vkqax6;
assign vis_r2_o[1] = Vmqax6;
assign vis_r2_o[25] = Uoqax6;
assign vis_r2_o[21] = Uqqax6;
assign vis_r2_o[20] = Usqax6;
assign vis_r2_o[19] = Uuqax6;
assign vis_r2_o[18] = Uwqax6;
assign vis_r2_o[17] = Uyqax6;
assign vis_r2_o[16] = U0rax6;
assign vis_r2_o[14] = U2rax6;
assign vis_r2_o[13] = U4rax6;
assign vis_r2_o[12] = U6rax6;
assign vis_r2_o[10] = U8rax6;
assign vis_r2_o[9] = Uarax6;
assign vis_r2_o[8] = Tcrax6;
assign vis_r8_o[2] = Serax6;
assign vis_r8_o[4] = Rgrax6;
assign vis_r8_o[23] = Qirax6;
assign vis_r8_o[30] = Qkrax6;
assign vis_r8_o[31] = Qmrax6;
assign vis_r8_o[0] = Qorax6;
assign vis_r8_o[1] = Pqrax6;
assign vis_r8_o[25] = Osrax6;
assign vis_r8_o[21] = Ourax6;
assign vis_r8_o[20] = Owrax6;
assign vis_r8_o[19] = Oyrax6;
assign vis_r8_o[18] = O0sax6;
assign vis_r8_o[17] = O2sax6;
assign vis_r8_o[16] = O4sax6;
assign vis_r8_o[14] = O6sax6;
assign vis_r8_o[13] = O8sax6;
assign vis_r8_o[12] = Oasax6;
assign vis_r8_o[10] = Ocsax6;
assign vis_r8_o[9] = Oesax6;
assign vis_r8_o[8] = Ngsax6;
assign vis_r12_o[2] = Misax6;
assign vis_r12_o[4] = Lksax6;
assign vis_r12_o[23] = Kmsax6;
assign vis_r12_o[30] = Kosax6;
assign vis_r12_o[31] = Kqsax6;
assign vis_r12_o[0] = Kssax6;
assign vis_r12_o[3] = Jusax6;
assign vis_r12_o[5] = Iwsax6;
assign vis_r12_o[6] = Hysax6;
assign vis_r12_o[7] = G0tax6;
assign vis_r12_o[24] = F2tax6;
assign vis_r12_o[26] = F4tax6;
assign vis_r12_o[27] = F6tax6;
assign vis_r12_o[29] = F8tax6;
assign vis_r12_o[1] = Fatax6;
assign vis_r12_o[25] = Ectax6;
assign vis_r12_o[21] = Eetax6;
assign vis_r12_o[20] = Egtax6;
assign vis_r12_o[19] = Eitax6;
assign vis_r12_o[18] = Ektax6;
assign vis_r12_o[17] = Emtax6;
assign vis_r12_o[16] = Eotax6;
assign vis_r12_o[14] = Eqtax6;
assign vis_r12_o[13] = Estax6;
assign vis_r12_o[12] = Eutax6;
assign vis_r12_o[10] = Ewtax6;
assign vis_r12_o[8] = Eytax6;
assign vis_r4_o[2] = D0uax6;
assign vis_r4_o[4] = C2uax6;
assign vis_r4_o[23] = B4uax6;
assign vis_r4_o[30] = B6uax6;
assign vis_r4_o[31] = B8uax6;
assign vis_r4_o[0] = Bauax6;
assign vis_r4_o[3] = Acuax6;
assign vis_r4_o[5] = Zduax6;
assign vis_r4_o[6] = Yfuax6;
assign vis_r4_o[7] = Xhuax6;
assign vis_r4_o[24] = Wjuax6;
assign vis_r4_o[26] = Wluax6;
assign vis_r4_o[27] = Wnuax6;
assign vis_r4_o[29] = Wpuax6;
assign vis_r4_o[1] = Wruax6;
assign vis_r4_o[25] = Vtuax6;
assign vis_r4_o[21] = Vvuax6;
assign vis_r4_o[20] = Vxuax6;
assign vis_r4_o[19] = Vzuax6;
assign vis_r4_o[18] = V1vax6;
assign vis_r4_o[17] = V3vax6;
assign vis_r4_o[16] = V5vax6;
assign vis_r4_o[14] = V7vax6;
assign vis_r4_o[13] = V9vax6;
assign vis_r4_o[12] = Vbvax6;
assign vis_r4_o[10] = Vdvax6;
assign vis_r4_o[9] = Vfvax6;
assign vis_r4_o[8] = Uhvax6;
assign vis_r7_o[2] = Tjvax6;
assign vis_r7_o[4] = Slvax6;
assign vis_r7_o[23] = Rnvax6;
assign vis_r7_o[30] = Rpvax6;
assign vis_r7_o[31] = Rrvax6;
assign vis_r7_o[0] = Rtvax6;
assign vis_r7_o[3] = Qvvax6;
assign vis_r7_o[5] = Pxvax6;
assign vis_r7_o[6] = Ozvax6;
assign vis_r7_o[7] = N1wax6;
assign vis_r7_o[24] = M3wax6;
assign vis_r7_o[26] = M5wax6;
assign vis_r7_o[27] = M7wax6;
assign vis_r7_o[29] = M9wax6;
assign vis_r7_o[1] = Mbwax6;
assign vis_r7_o[25] = Ldwax6;
assign vis_r7_o[21] = Lfwax6;
assign vis_r7_o[20] = Lhwax6;
assign vis_r7_o[19] = Ljwax6;
assign vis_r7_o[18] = Llwax6;
assign vis_r7_o[17] = Lnwax6;
assign vis_r7_o[16] = Lpwax6;
assign vis_r7_o[14] = Lrwax6;
assign vis_r7_o[13] = Ltwax6;
assign vis_r7_o[12] = Lvwax6;
assign vis_r7_o[10] = Lxwax6;
assign vis_r7_o[8] = Lzwax6;
assign vis_r3_o[2] = K1xax6;
assign vis_r3_o[4] = J3xax6;
assign Jfgpw6[1] = I5xax6;
assign Bagpw6[23] = J7xax6;
assign Bagpw6[15] = L9xax6;
assign Tzfpw6[15] = Nbxax6;
assign Bagpw6[14] = Pdxax6;
assign Tzfpw6[14] = Rfxax6;
assign Bagpw6[7] = Thxax6;
assign Tzfpw6[7] = Ujxax6;
assign Bagpw6[2] = Vlxax6;
assign Bagpw6[1] = Wnxax6;
assign Fkfpw6[13] = Xpxax6;
assign Fkfpw6[2] = Xrxax6;
assign Fkfpw6[4] = Wtxax6;
assign vis_r3_o[23] = Vvxax6;
assign vis_r3_o[30] = Vxxax6;
assign vis_r3_o[31] = Vzxax6;
assign vis_r3_o[0] = V1yax6;
assign vis_r3_o[3] = U3yax6;
assign Fkfpw6[3] = T5yax6;
assign vis_r3_o[5] = S7yax6;
assign Jfgpw6[3] = R9yax6;
assign Evdpw6 = (!Sbyax6);
assign Ahghu6 = Pdyax6;
assign R4gpw6[41] = Mfyax6;
assign R4gpw6[42] = Ohyax6;
assign R4gpw6[43] = Qjyax6;
assign R4gpw6[45] = Slyax6;
assign R4gpw6[46] = Unyax6;
assign R4gpw6[47] = Wpyax6;
assign R4gpw6[11] = Yryax6;
assign R4gpw6[13] = Auyax6;
assign R4gpw6[14] = Cwyax6;
assign R4gpw6[15] = Eyyax6;
assign Qqdhu6 = G0zax6;
assign Ndghu6 = I2zax6;
assign R4gpw6[33] = H4zax6;
assign R4gpw6[34] = J6zax6;
assign R4gpw6[35] = L8zax6;
assign R4gpw6[37] = Nazax6;
assign R4gpw6[38] = Pczax6;
assign R4gpw6[39] = Rezax6;
assign R4gpw6[7] = Tgzax6;
assign R4gpw6[6] = Uizax6;
assign R4gpw6[5] = Vkzax6;
assign R4gpw6[3] = Wmzax6;
assign R4gpw6[2] = Xozax6;
assign R4gpw6[1] = Yqzax6;
assign Bxghu6 = Zszax6;
assign Dvghu6 = Avzax6;
assign Vbgpw6[1] = Cxzax6;
assign Vbgpw6[5] = Czzax6;
assign Vbgpw6[7] = C10bx6;
assign Vbgpw6[8] = C30bx6;
assign Vbgpw6[10] = C50bx6;
assign Vbgpw6[11] = D70bx6;
assign Vbgpw6[12] = E90bx6;
assign Vbgpw6[13] = Fb0bx6;
assign Vbgpw6[14] = Gd0bx6;
assign Vbgpw6[15] = Hf0bx6;
assign Vbgpw6[16] = Ih0bx6;
assign Vbgpw6[17] = Jj0bx6;
assign Vbgpw6[18] = Kl0bx6;
assign Vbgpw6[19] = Ln0bx6;
assign Vbgpw6[20] = Mp0bx6;
assign Vbgpw6[21] = Nr0bx6;
assign Vbgpw6[23] = Ot0bx6;
assign Vbgpw6[25] = Pv0bx6;
assign Vbgpw6[27] = Qx0bx6;
assign Vbgpw6[30] = Rz0bx6;
assign Xudpw6 = (!S11bx6);
assign Odgpw6[0] = U31bx6;
assign Qudpw6 = (!W51bx6);
assign Odgpw6[12] = Z71bx6;
assign Judpw6 = (!Ca1bx6);
assign Odgpw6[10] = Fc1bx6;
assign Cudpw6 = (!Ie1bx6);
assign Odgpw6[11] = Lg1bx6;
assign Vtdpw6 = (!Oi1bx6);
assign Odgpw6[13] = Rk1bx6;
assign Otdpw6 = (!Um1bx6);
assign Odgpw6[14] = Xo1bx6;
assign Htdpw6 = (!Ar1bx6);
assign Odgpw6[17] = Dt1bx6;
assign Atdpw6 = (!Gv1bx6);
assign Odgpw6[16] = Jx1bx6;
assign Tsdpw6 = (!Mz1bx6);
assign Odgpw6[18] = P12bx6;
assign Msdpw6 = (!S32bx6);
assign Odgpw6[19] = V52bx6;
assign Fsdpw6 = (!Y72bx6);
assign Odgpw6[1] = Aa2bx6;
assign Yrdpw6 = (!Cc2bx6);
assign Odgpw6[20] = Fe2bx6;
assign Rrdpw6 = (!Ig2bx6);
assign Odgpw6[21] = Li2bx6;
assign Krdpw6 = (!Ok2bx6);
assign Odgpw6[25] = Rm2bx6;
assign Drdpw6 = (!Uo2bx6);
assign Odgpw6[23] = Xq2bx6;
assign Wqdpw6 = (!At2bx6);
assign Odgpw6[24] = Dv2bx6;
assign Pqdpw6 = (!Gx2bx6);
assign Odgpw6[26] = Jz2bx6;
assign Iqdpw6 = (!M13bx6);
assign Odgpw6[27] = P33bx6;
assign Bqdpw6 = (!S53bx6);
assign Odgpw6[28] = V73bx6;
assign Updpw6 = (!Y93bx6);
assign Odgpw6[29] = Bc3bx6;
assign Npdpw6 = (!Ee3bx6);
assign Odgpw6[31] = Hg3bx6;
assign Gpdpw6 = (!Ki3bx6);
assign Odgpw6[5] = Mk3bx6;
assign Zodpw6 = (!Om3bx6);
assign Odgpw6[7] = Qo3bx6;
assign Sodpw6 = (!Sq3bx6);
assign Odgpw6[8] = Us3bx6;
assign R4gpw6[49] = Wu3bx6;
assign R4gpw6[50] = Yw3bx6;
assign R4gpw6[51] = Az3bx6;
assign R4gpw6[53] = C14bx6;
assign R4gpw6[54] = E34bx6;
assign R4gpw6[55] = G54bx6;
assign R4gpw6[17] = I74bx6;
assign R4gpw6[18] = K94bx6;
assign R4gpw6[19] = Mb4bx6;
assign R4gpw6[21] = Od4bx6;
assign R4gpw6[22] = Qf4bx6;
assign R4gpw6[23] = Sh4bx6;
assign B3gpw6[1] = Uj4bx6;
assign B3gpw6[0] = Tl4bx6;
assign R4gpw6[57] = Sn4bx6;
assign R4gpw6[58] = Up4bx6;
assign R4gpw6[59] = Wr4bx6;
assign R4gpw6[61] = Yt4bx6;
assign R4gpw6[62] = Aw4bx6;
assign R4gpw6[63] = Cy4bx6;
assign R4gpw6[25] = E05bx6;
assign R4gpw6[26] = G25bx6;
assign R4gpw6[27] = I45bx6;
assign R4gpw6[29] = K65bx6;
assign R4gpw6[30] = M85bx6;
assign R4gpw6[31] = Oa5bx6;
assign Fkfpw6[5] = Qc5bx6;
assign vis_r3_o[6] = Pe5bx6;
assign vis_r3_o[7] = Og5bx6;
assign vis_r3_o[24] = Ni5bx6;
assign vis_r3_o[26] = Nk5bx6;
assign vis_r3_o[27] = Nm5bx6;
assign vis_r3_o[29] = No5bx6;
assign vis_r3_o[1] = Nq5bx6;
assign Iwfpw6[1] = Ms5bx6;
assign Fkfpw6[1] = Nu5bx6;
assign vis_pc_o[10] = Mw5bx6;
assign vis_r3_o[25] = Jy5bx6;
assign vis_pc_o[8] = J06bx6;
assign L8ehu6 = F26bx6;
assign vis_r3_o[21] = D46bx6;
assign vis_r3_o[20] = D66bx6;
assign vis_r3_o[19] = D86bx6;
assign vis_r3_o[18] = Da6bx6;
assign vis_r3_o[17] = Dc6bx6;
assign vis_r3_o[16] = De6bx6;
assign vis_r3_o[14] = Dg6bx6;
assign vis_r3_o[13] = Di6bx6;
assign vis_r3_o[12] = Dk6bx6;
assign Fkfpw6[12] = Dm6bx6;
assign vis_r3_o[10] = Do6bx6;
assign vis_r3_o[9] = Dq6bx6;
assign vis_r3_o[8] = Cs6bx6;
assign Uthpw6[11] = Bu6bx6;
assign Iahpw6[10] = Gw6bx6;
assign Shhpw6[11] = Xx6bx6;
assign Fkfpw6[11] = C07bx6;
assign vis_r0_o[11] = C27bx6;
assign vis_r1_o[11] = C47bx6;
assign vis_r2_o[11] = C67bx6;
assign vis_r3_o[11] = C87bx6;
assign vis_r8_o[11] = Ca7bx6;
assign vis_r9_o[11] = Cc7bx6;
assign vis_r10_o[11] = Ce7bx6;
assign vis_r11_o[11] = Cg7bx6;
assign vis_r4_o[11] = Ci7bx6;
assign vis_r5_o[11] = Ck7bx6;
assign vis_r6_o[11] = Cm7bx6;
assign vis_r7_o[11] = Co7bx6;
assign vis_pc_o[14] = Cq7bx6;
assign vis_r0_o[15] = Zr7bx6;
assign vis_r1_o[15] = Zt7bx6;
assign vis_r2_o[15] = Zv7bx6;
assign vis_r3_o[15] = Zx7bx6;
assign vis_r8_o[15] = Zz7bx6;
assign vis_r9_o[15] = Z18bx6;
assign vis_r10_o[15] = Z38bx6;
assign vis_r11_o[15] = Z58bx6;
assign vis_r4_o[15] = Z78bx6;
assign vis_r5_o[15] = Z98bx6;
assign vis_r6_o[15] = Zb8bx6;
assign vis_r7_o[15] = Zd8bx6;
assign vis_r12_o[15] = Zf8bx6;
assign vis_r14_o[15] = Zh8bx6;
assign vis_msp_o[13] = Zj8bx6;
assign vis_psp_o[13] = Zl8bx6;
assign vis_r12_o[11] = Zn8bx6;
assign vis_r14_o[11] = Zp8bx6;
assign vis_msp_o[9] = Zr8bx6;
assign vis_psp_o[9] = Yt8bx6;
assign K7hpw6[11] = Xv8bx6;
assign E1hpw6[11] = Ux8bx6;
assign Gtgpw6[11] = Rz8bx6;
assign Trgpw6[11] = N19bx6;
assign Gqgpw6[11] = J39bx6;
assign Togpw6[11] = F59bx6;
assign Jshpw6[11] = B79bx6;
assign Shhpw6[6] = Q89bx6;
assign Fkfpw6[6] = Ua9bx6;
assign K7hpw6[6] = Tc9bx6;
assign E1hpw6[6] = Pe9bx6;
assign Gtgpw6[6] = Lg9bx6;
assign Trgpw6[6] = Hi9bx6;
assign Gqgpw6[6] = Dk9bx6;
assign Togpw6[6] = Zl9bx6;
assign Jshpw6[6] = Vn9bx6;
assign Lodpw6 = (!Jp9bx6);
assign Odgpw6[6] = Lr9bx6;
assign Vbgpw6[6] = Nt9bx6;
assign R4gpw6[0] = Nv9bx6;
assign Bagpw6[6] = Ox9bx6;
assign R4gpw6[56] = Pz9bx6;
assign R4gpw6[48] = R1abx6;
assign R4gpw6[40] = T3abx6;
assign R4gpw6[32] = V5abx6;
assign R4gpw6[24] = X7abx6;
assign R4gpw6[16] = Z9abx6;
assign R4gpw6[8] = Bcabx6;
assign Uthpw6[5] = Ceabx6;
assign Uthpw6[13] = Ggabx6;
assign Shhpw6[14] = Liabx6;
assign K7hpw6[14] = Qkabx6;
assign E1hpw6[14] = Nmabx6;
assign Gtgpw6[14] = Koabx6;
assign Trgpw6[14] = Hqabx6;
assign Gqgpw6[14] = Esabx6;
assign Togpw6[14] = Buabx6;
assign Jshpw6[14] = Yvabx6;
assign vis_pc_o[21] = Nxabx6;
assign Tzfpw6[2] = Kzabx6;
assign Vbgpw6[2] = L1bbx6;
assign Eodpw6 = (!L3bbx6);
assign Odgpw6[2] = N5bbx6;
assign vis_pc_o[9] = P7bbx6;
assign Uthpw6[1] = L9bbx6;
assign Fkfpw6[17] = Pbbbx6;
assign Uthpw6[17] = Pdbbx6;
assign Iahpw6[16] = Ufbbx6;
assign Shhpw6[17] = Lhbbx6;
assign K7hpw6[17] = Qjbbx6;
assign E1hpw6[17] = Nlbbx6;
assign Gtgpw6[17] = Knbbx6;
assign Trgpw6[17] = Hpbbx6;
assign Gqgpw6[17] = Erbbx6;
assign Togpw6[17] = Btbbx6;
assign Jshpw6[17] = Yubbx6;
assign Fkfpw6[25] = Nwbbx6;
assign Fkfpw6[27] = Nybbx6;
assign Uthpw6[27] = N0cbx6;
assign Iahpw6[26] = S2cbx6;
assign Iahpw6[25] = J4cbx6;
assign Shhpw6[26] = A6cbx6;
assign Fkfpw6[26] = F8cbx6;
assign K7hpw6[26] = Facbx6;
assign E1hpw6[26] = Cccbx6;
assign Gtgpw6[26] = Zdcbx6;
assign Trgpw6[26] = Wfcbx6;
assign Gqgpw6[26] = Thcbx6;
assign Togpw6[26] = Qjcbx6;
assign Jshpw6[26] = Nlcbx6;
assign Uthpw6[26] = Cncbx6;
assign Zbhpw6[26] = Hpcbx6;
assign Shhpw6[27] = Drcbx6;
assign K7hpw6[27] = Itcbx6;
assign E1hpw6[27] = Fvcbx6;
assign Gtgpw6[27] = Cxcbx6;
assign Trgpw6[27] = Zycbx6;
assign Gqgpw6[27] = W0dbx6;
assign Togpw6[27] = T2dbx6;
assign Jshpw6[27] = Q4dbx6;
assign Fkfpw6[30] = F6dbx6;
assign Uthpw6[23] = F8dbx6;
assign Iahpw6[22] = Kadbx6;
assign Iahpw6[21] = Bcdbx6;
assign Iahpw6[20] = Sddbx6;
assign Iahpw6[19] = Jfdbx6;
assign Shhpw6[20] = Ahdbx6;
assign Fkfpw6[20] = Fjdbx6;
assign K7hpw6[20] = Fldbx6;
assign E1hpw6[20] = Cndbx6;
assign Gtgpw6[20] = Zodbx6;
assign Trgpw6[20] = Wqdbx6;
assign Gqgpw6[20] = Tsdbx6;
assign Togpw6[20] = Qudbx6;
assign Jshpw6[20] = Nwdbx6;
assign Uthpw6[20] = Cydbx6;
assign Shhpw6[21] = H0ebx6;
assign Fkfpw6[21] = M2ebx6;
assign K7hpw6[21] = M4ebx6;
assign E1hpw6[21] = J6ebx6;
assign Gtgpw6[21] = G8ebx6;
assign Trgpw6[21] = Daebx6;
assign Gqgpw6[21] = Acebx6;
assign Togpw6[21] = Xdebx6;
assign Jshpw6[21] = Ufebx6;
assign Uthpw6[21] = Jhebx6;
assign Shhpw6[22] = Ojebx6;
assign Fkfpw6[22] = Tlebx6;
assign vis_r0_o[22] = Tnebx6;
assign vis_r1_o[22] = Tpebx6;
assign vis_r2_o[22] = Trebx6;
assign vis_r3_o[22] = Ttebx6;
assign vis_r8_o[22] = Tvebx6;
assign vis_r9_o[22] = Txebx6;
assign vis_r10_o[22] = Tzebx6;
assign vis_r11_o[22] = T1fbx6;
assign vis_r4_o[22] = T3fbx6;
assign vis_r5_o[22] = T5fbx6;
assign vis_r6_o[22] = T7fbx6;
assign vis_r7_o[22] = T9fbx6;
assign vis_r12_o[22] = Tbfbx6;
assign vis_r14_o[22] = Tdfbx6;
assign vis_msp_o[20] = Tffbx6;
assign vis_psp_o[20] = Thfbx6;
assign K7hpw6[22] = Tjfbx6;
assign E1hpw6[22] = Qlfbx6;
assign Gtgpw6[22] = Nnfbx6;
assign Trgpw6[22] = Kpfbx6;
assign Gqgpw6[22] = Hrfbx6;
assign Togpw6[22] = Etfbx6;
assign Jshpw6[22] = Bvfbx6;
assign Uthpw6[22] = Qwfbx6;
assign Xndpw6 = (!Vyfbx6);
assign Odgpw6[22] = Y0gbx6;
assign Vbgpw6[22] = B3gbx6;
assign R4gpw6[4] = C5gbx6;
assign Bagpw6[22] = D7gbx6;
assign Tzfpw6[22] = F9gbx6;
assign R4gpw6[60] = Hbgbx6;
assign R4gpw6[52] = Jdgbx6;
assign R4gpw6[44] = Lfgbx6;
assign R4gpw6[36] = Nhgbx6;
assign R4gpw6[28] = Pjgbx6;
assign R4gpw6[20] = Rlgbx6;
assign R4gpw6[12] = Tngbx6;
assign L1gpw6[0] = Vpgbx6;
assign Shhpw6[23] = Urgbx6;
assign Fkfpw6[23] = Ztgbx6;
assign K7hpw6[23] = Zvgbx6;
assign E1hpw6[23] = Wxgbx6;
assign Gtgpw6[23] = Tzgbx6;
assign Trgpw6[23] = Q1hbx6;
assign Gqgpw6[23] = N3hbx6;
assign Togpw6[23] = K5hbx6;
assign Jshpw6[23] = H7hbx6;
assign Ppfpw6[15] = W8hbx6;
assign K7hpw6[29] = Wahbx6;
assign E1hpw6[29] = Tchbx6;
assign Tnhpw6[0] = Qehbx6;
assign Qndpw6 = (!Eghbx6);
assign Odgpw6[4] = Gihbx6;
assign Vbgpw6[4] = Ikhbx6;
assign Bagpw6[4] = Imhbx6;
assign Tzfpw6[4] = Johbx6;
assign Gfghu6 = Kqhbx6;
assign Jndpw6 = (!Kshbx6);
assign Odgpw6[3] = Muhbx6;
assign Vbgpw6[3] = Owhbx6;
assign Bagpw6[3] = Oyhbx6;
assign Tzfpw6[3] = P0ibx6;
assign Jshpw6[25] = Q2ibx6;
assign Vxmhu6 = F4ibx6;
assign vis_apsr_o[0] = X5ibx6;
assign vis_r2_o[28] = R7ibx6;
assign vis_r3_o[28] = R9ibx6;
assign vis_r8_o[28] = Rbibx6;
assign vis_r9_o[28] = Rdibx6;
assign vis_r10_o[28] = Rfibx6;
assign vis_r4_o[28] = Rhibx6;
assign vis_r5_o[28] = Rjibx6;
assign vis_r6_o[28] = Rlibx6;
assign vis_r7_o[28] = Rnibx6;
assign vis_r12_o[28] = Rpibx6;
assign vis_r14_o[28] = Rribx6;
assign vis_psp_o[26] = Rtibx6;
assign vis_r12_o[9] = Rvibx6;
assign vis_r14_o[9] = Qxibx6;
assign vis_msp_o[7] = Pzibx6;
assign vis_psp_o[7] = O1jbx6;
assign K7hpw6[9] = N3jbx6;
assign E1hpw6[9] = J5jbx6;
assign Gtgpw6[9] = F7jbx6;
assign Trgpw6[9] = B9jbx6;
assign Gqgpw6[9] = Xajbx6;
assign Togpw6[9] = Tcjbx6;
assign vis_msp_o[26] = Pejbx6;
assign Cndpw6 = (!Pgjbx6);
assign Odgpw6[9] = Rijbx6;
assign Vbgpw6[9] = Tkjbx6;
assign Bagpw6[9] = Tmjbx6;
assign Tzfpw6[9] = Uojbx6;
assign Hrfpw6[3] = Vqjbx6;
assign Hrfpw6[2] = Usjbx6;
assign Hrfpw6[1] = Tujbx6;
assign Hrfpw6[14] = Swjbx6;
assign Fkfpw6[18] = Syjbx6;
assign Vbgpw6[31] = S0kbx6;
assign Krghu6 = T2kbx6;
assign Iwfpw6[0] = S4kbx6;
assign Fkfpw6[19] = T6kbx6;
assign Righu6 = T8kbx6;
assign Jydhu6 = Qakbx6;
assign Uthpw6[7] = Nckbx6;
assign SYSRESETREQ = Rekbx6;
assign Kaohu6 = (!Rekbx6);
assign Fkfpw6[24] = Tgkbx6;
assign Aygpw6[0] = Tikbx6;
assign G4hpw6[0] = Pkkbx6;
assign Dhgpw6[0] = Lmkbx6;
assign Qnghu6 = Cokbx6;
assign SWDOEN = Dqkbx6;
assign Vrkbx6 = ({{Jshpw6[9:4], Tnhpw6}, 1'b0} + {{1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, Aphpw6, E4yhu6}, 1'b1});
assign Gmhpw6 = Vrkbx6[33:1];
assign Yuhhu6 = (({R9ohu6, Mzihu6, Eyihu6, Wwihu6, Ovihu6, Guihu6,
 Ysihu6, Qrihu6, Iqihu6, Apihu6, Snihu6, Kmihu6, Clihu6, Ujihu6,
 Miihu6, Ehihu6, Wfihu6, Oeihu6, Gdihu6, Ybihu6, Qaihu6, I9ihu6,
 A8ihu6, S6ihu6, K5ihu6, C4ihu6, U2ihu6, M1ihu6, E0ihu6, Wyhhu6,
 Oxhhu6, Gwhhu6} == {E1hpw6, Edkhu6, Wbkhu6}) ? 1'b1 : 1'b0);
assign Ntkbx6 = ({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
 1'b1, 1'b1, 1'b1} << {Oakhu6, G9khu6, Y7khu6, Q6khu6, I5khu6});
assign {K5epw6, U0jhu6, C2jhu6, K3jhu6, S4jhu6, A6jhu6, I7jhu6, Q8jhu6,
 Y9jhu6, Gbjhu6, Ocjhu6, Wdjhu6, Efjhu6, Mgjhu6, Uhjhu6, Cjjhu6,
 Kkjhu6, Sljhu6, Anjhu6, Iojhu6, Qpjhu6, Yqjhu6, Gsjhu6, Otjhu6,
 Wujhu6, Ewjhu6, Mxjhu6, Uyjhu6, C0khu6, K1khu6, S2khu6, A4khu6}
 = Ntkbx6[31:0];
assign Mekhu6 = (({M9ohu6, Uilhu6, Nhlhu6, Gglhu6, Zelhu6, Sdlhu6,
 Lclhu6, Eblhu6, W9lhu6, O8lhu6, G7lhu6, Y5lhu6, Q4lhu6, I3lhu6,
 A2lhu6, S0lhu6, Kzkhu6, Cykhu6, Uwkhu6, Mvkhu6, Eukhu6, Wskhu6,
 Orkhu6, Gqkhu6, Yokhu6, Qnkhu6, Imkhu6, Alkhu6, Sjkhu6, Kikhu6,
 Chkhu6, Ufkhu6} == {K7hpw6, Avmhu6, Ttmhu6}) ? 1'b1 : 1'b0);
assign Nvkbx6 = ({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
 1'b1, 1'b1, 1'b1} << {Msmhu6, Frmhu6, Ypmhu6, Romhu6, Knmhu6});
assign {H6epw6, Bklhu6, Illhu6, Pmlhu6, Wnlhu6, Dplhu6, Kqlhu6, Rrlhu6,
 Yslhu6, Fulhu6, Mvlhu6, Twlhu6, Aylhu6, Hzlhu6, O0mhu6, V1mhu6,
 C3mhu6, J4mhu6, Q5mhu6, X6mhu6, E8mhu6, L9mhu6, Samhu6, Zbmhu6,
 Gdmhu6, Nemhu6, Ufmhu6, Bhmhu6, Iimhu6, Pjmhu6, Wkmhu6, Dmmhu6}
 = Nvkbx6[31:0];
assign Wphhu6 = (({V0epw6, O0epw6, H0epw6, A0epw6, Tzdpw6, Mzdpw6,
 Fzdpw6, Yydpw6, Rydpw6, Kydpw6, Dydpw6, Wxdpw6, Pxdpw6,
 Tugpw6[13:11], Ixdpw6, Tugpw6[9:0]} == Togpw6) ? 1'b1 : 1'b0);
assign Drhhu6 = (({V0epw6, O0epw6, H0epw6, A0epw6, Tzdpw6, Mzdpw6,
 Fzdpw6, Yydpw6, Rydpw6, Kydpw6, Dydpw6, Wxdpw6, Pxdpw6,
 Tugpw6[13:11], Ixdpw6, Tugpw6[9:0]} == Gqgpw6) ? 1'b1 : 1'b0);
assign Kshhu6 = (({V0epw6, O0epw6, H0epw6, A0epw6, Tzdpw6, Mzdpw6,
 Fzdpw6, Yydpw6, Rydpw6, Kydpw6, Dydpw6, Wxdpw6, Pxdpw6,
 Tugpw6[13:11], Ixdpw6, Tugpw6[9:0]} == Trgpw6) ? 1'b1 : 1'b0);
assign Rthhu6 = (({V0epw6, O0epw6, H0epw6, A0epw6, Tzdpw6, Mzdpw6,
 Fzdpw6, Yydpw6, Rydpw6, Kydpw6, Dydpw6, Wxdpw6, Pxdpw6,
 Tugpw6[13:11], Ixdpw6, Tugpw6[9:0]} == Gtgpw6) ? 1'b1 : 1'b0);
assign L6gpw6 = (Tzfpw6 - 1'b1);
assign {Xlfpw6, E7epw6} = ({Vnfpw6, X5phu6} - 1'b1);
assign Zsfpw6 = (vis_pc_o + 1'b1);
assign {N5fpw6, B8epw6} = ({vis_pc_o[30:2], R0ghu6} + 1'b1);
assign {Y8epw6, V9epw6, Saepw6, Pbepw6, Mcepw6, Jdepw6, Heepw6, Ffepw6,
 Dgepw6, Bhepw6, Zhepw6, Xiepw6, Vjepw6, Tkepw6, Rlepw6, Pmepw6,
 Nnepw6, Loepw6, Jpepw6, Hqepw6, Frepw6, Dsepw6, Btepw6, Ztepw6,
 Xuepw6, Vvepw6, Twepw6, Rxepw6, Pyepw6, Nzepw6, L0fpw6, J1fpw6,
 Affpw6} = (Mifpw6 * Tgfpw6);
assign Nxkbx6 = ({{Qbehu6, Edehu6, Seehu6, Ggehu6, Uhehu6, Ijehu6,
 Wkehu6, Kmehu6, Ynehu6, Mpehu6, Arehu6, Osehu6, Cuehu6, Qvehu6,
 Exehu6, Syehu6, G0fhu6, U1fhu6, I3fhu6, W4fhu6, K6fhu6, Y7fhu6,
 M9fhu6, Abfhu6, Ocfhu6, Cefhu6, Qffhu6, Dhfhu6, Qifhu6, Dkfhu6,
 Qlfhu6, Dnfhu6, Qofhu6}, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Dqfhu6}, 1'b1});
assign {Caehu6, Eafpw6} = Nxkbx6[33:1];
assign Ozkbx6 = ({{1'b0, Idfpw6}, 1'b0} + {{1'b0, D5epw6, Qbfpw6[30:23],
 P4epw6, I4epw6, B4epw6, U3epw6, N3epw6, G3epw6, Z2epw6, L2epw6,
 X1epw6, Q1epw6, J1epw6, C1epw6, Qbfpw6[10], Q5phu6, W4epw6,
 S2epw6, E2epw6, Qbfpw6[5:0]}, 1'b1});
assign {Qbehu6, Edehu6, Seehu6, Ggehu6, Uhehu6, Ijehu6, Wkehu6, Kmehu6,
 Ynehu6, Mpehu6, Arehu6, Osehu6, Cuehu6, Qvehu6, Exehu6, Syehu6,
 G0fhu6, U1fhu6, I3fhu6, W4fhu6, K6fhu6, Y7fhu6, M9fhu6, Abfhu6,
 Ocfhu6, Cefhu6, Qffhu6, Dhfhu6, Qifhu6, Dkfhu6, Qlfhu6, Dnfhu6,
 Qofhu6} = Ozkbx6[33:1];
assign I5nhu6 = (~(L4yhu6 & S4yhu6));
assign S4yhu6 = (~(Z4yhu6 & SWDOEN));
assign L4yhu6 = (G5yhu6 & N5yhu6);
assign G5yhu6 = (~(U5yhu6 & B6yhu6));
assign B6yhu6 = (~(I6yhu6 & P6yhu6));
assign P6yhu6 = (~(W6yhu6 & D7yhu6));
assign D7yhu6 = (~(K7yhu6 | Ighpw6[4]));
assign W6yhu6 = (~(R7yhu6 | Y7yhu6));
assign Zehpw6[6] = (~(F8yhu6 & M8yhu6));
assign M8yhu6 = (~(T8yhu6 & Fnnhu6));
assign F8yhu6 = (A9yhu6 & H9yhu6);
assign H9yhu6 = (~(O9yhu6 & V9yhu6));
assign V9yhu6 = (~(Cayhu6 & Jayhu6));
assign A9yhu6 = (~(U5yhu6 & Qayhu6));
assign Qayhu6 = (~(Xayhu6 & Ebyhu6));
assign Ebyhu6 = (~(Lbyhu6 | Sbyhu6));
assign Xayhu6 = (Zbyhu6 & Gcyhu6);
assign Gcyhu6 = (~(Ighpw6[4] & Ncyhu6));
assign Ncyhu6 = (~(Ucyhu6 & Bdyhu6));
assign Bdyhu6 = (Ighpw6[1] | Ighpw6[2]);
assign Ucyhu6 = (Idyhu6 & Pdyhu6);
assign Idyhu6 = (Wdyhu6 | Deyhu6);
assign Zbyhu6 = (Mdhpw6[3] ? Reyhu6 : Keyhu6);
assign Reyhu6 = (Yeyhu6 & Ffyhu6);
assign Yeyhu6 = (Mfyhu6 & Tfyhu6);
assign Keyhu6 = (~(Agyhu6 | Hgyhu6));
assign Zehpw6[5] = (~(Ogyhu6 & Vgyhu6));
assign Vgyhu6 = (~(O9yhu6 & Mdhpw6[3]));
assign Ogyhu6 = (Chyhu6 & Jhyhu6);
assign Jhyhu6 = (~(Qhyhu6 & U5yhu6));
assign Qhyhu6 = (Xhyhu6 & Eiyhu6);
assign Xhyhu6 = (~(Liyhu6 & Siyhu6));
assign Siyhu6 = (~(Ziyhu6 & Mdhpw6[0]));
assign Liyhu6 = (~(Ighpw6[2] & Gjyhu6));
assign Chyhu6 = (~(T8yhu6 & Njyhu6));
assign Njyhu6 = (~(Ujyhu6 ^ Bkyhu6));
assign Bkyhu6 = (Ikyhu6 & Pkyhu6);
assign Ikyhu6 = (~(Eiyhu6 | Wdyhu6));
assign Zehpw6[4] = (~(Wkyhu6 & Dlyhu6));
assign Dlyhu6 = (Klyhu6 & Rlyhu6);
assign Klyhu6 = (~(Ylyhu6 & Fmyhu6));
assign Ylyhu6 = (~(Mmyhu6 | B7nhu6));
assign Wkyhu6 = (Tmyhu6 & Anyhu6);
assign Anyhu6 = (~(U5yhu6 & Hnyhu6));
assign Hnyhu6 = (Onyhu6 | Vnyhu6);
assign Onyhu6 = (~(Coyhu6 & Joyhu6));
assign Coyhu6 = (Eiyhu6 | I6yhu6);
assign Tmyhu6 = (~(T8yhu6 & Qoyhu6));
assign Qoyhu6 = (Xoyhu6 | Epyhu6);
assign Xoyhu6 = (Pkyhu6 ? Lpyhu6 : Ighpw6[4]);
assign Lpyhu6 = (~(Wdyhu6 | Ighpw6[4]));
assign Zehpw6[3] = (~(Spyhu6 & Zpyhu6));
assign Zpyhu6 = (~(U5yhu6 & Gqyhu6));
assign Gqyhu6 = (~(Nqyhu6 & Uqyhu6));
assign Uqyhu6 = (Bryhu6 & Iryhu6);
assign Bryhu6 = (Ffyhu6 | Mdhpw6[3]);
assign Ffyhu6 = (Pryhu6 & Wryhu6);
assign Nqyhu6 = (~(Dsyhu6 | Ksyhu6));
assign Dsyhu6 = (Ighpw6[3] ? Ysyhu6 : Rsyhu6);
assign Ysyhu6 = (!Ftyhu6);
assign Rsyhu6 = (~(Pdyhu6 | Ighpw6[4]));
assign Spyhu6 = (Mtyhu6 & N5yhu6);
assign Mtyhu6 = (~(T8yhu6 & Ttyhu6));
assign Ttyhu6 = (~(Wdyhu6 ^ Pkyhu6));
assign Zehpw6[2] = (~(Auyhu6 & Huyhu6));
assign Huyhu6 = (~(T8yhu6 & Ouyhu6));
assign Ouyhu6 = (~(Vuyhu6 ^ Cvyhu6));
assign Auyhu6 = (~(U5yhu6 & Jvyhu6));
assign Jvyhu6 = (~(Qvyhu6 & Xvyhu6));
assign Xvyhu6 = (Ewyhu6 & Lwyhu6);
assign Lwyhu6 = (~(Swyhu6 & Zwyhu6));
assign Ewyhu6 = (Gxyhu6 & Ftyhu6);
assign Gxyhu6 = (~(Mdhpw6[3] & Nxyhu6));
assign Nxyhu6 = (~(Uxyhu6 & Byyhu6));
assign Byyhu6 = (~(Iyyhu6 & Cvyhu6));
assign Uxyhu6 = (~(Pyyhu6 & Wyyhu6));
assign Wyyhu6 = (~(Dzyhu6 & Kzyhu6));
assign Kzyhu6 = (~(Lbyhu6 & Mdhpw6[0]));
assign Dzyhu6 = (Pryhu6 | Rzyhu6);
assign Qvyhu6 = (~(Ksyhu6 | Vnyhu6));
assign Vnyhu6 = (Mdhpw6[3] ? Hgyhu6 : Yzyhu6);
assign Yzyhu6 = (~(Mfyhu6 & Tfyhu6));
assign Ksyhu6 = (~(I6yhu6 & F0zhu6));
assign F0zhu6 = (~(M0zhu6 & Ziyhu6));
assign M0zhu6 = (~(Mdhpw6[0] | Ighpw6[4]));
assign I6yhu6 = (~(T0zhu6 | A1zhu6));
assign Zehpw6[1] = (~(H1zhu6 & O1zhu6));
assign O1zhu6 = (~(U5yhu6 & V1zhu6));
assign V1zhu6 = (~(C2zhu6 & J2zhu6));
assign J2zhu6 = (Q2zhu6 & X2zhu6);
assign X2zhu6 = (~(E3zhu6 & Ighpw6[0]));
assign E3zhu6 = (L3zhu6 & Eiyhu6);
assign L3zhu6 = (~(S3zhu6 & Z3zhu6));
assign Z3zhu6 = (Y7yhu6 | Mdhpw6[0]);
assign S3zhu6 = (Ighpw6[1] | Ighpw6[3]);
assign Q2zhu6 = (G4zhu6 & Joyhu6);
assign G4zhu6 = (~(N4zhu6 & U4zhu6));
assign N4zhu6 = (Hknhu6 & B5zhu6);
assign B5zhu6 = (~(Pyyhu6 & I5zhu6));
assign I5zhu6 = (P5zhu6 | R7yhu6);
assign C2zhu6 = (W5zhu6 & D6zhu6);
assign D6zhu6 = (Mdhpw6[3] ? R6zhu6 : K6zhu6);
assign R6zhu6 = (Mfyhu6 & Y6zhu6);
assign Y6zhu6 = (~(F7zhu6 & Lbyhu6));
assign Lbyhu6 = (M7zhu6 & T7zhu6);
assign F7zhu6 = (Mdhpw6[2] & A8zhu6);
assign A8zhu6 = (~(H8zhu6 & Mdhpw6[0]));
assign H8zhu6 = (~(O8zhu6 | Ulnhu6));
assign Mfyhu6 = (~(V8zhu6 & Epyhu6));
assign V8zhu6 = (~(C9zhu6 | Ighpw6[2]));
assign K6zhu6 = (Pryhu6 & Tfyhu6);
assign W5zhu6 = (J9zhu6 & Q9zhu6);
assign Q9zhu6 = (~(X9zhu6 & R7yhu6));
assign H1zhu6 = (Eazhu6 & Rlyhu6);
assign Rlyhu6 = (~(O9yhu6 & Cayhu6));
assign Eazhu6 = (~(T8yhu6 & Lazhu6));
assign Lazhu6 = (~(Deyhu6 & Sazhu6));
assign Sazhu6 = (Zazhu6 | Ighpw6[1]);
assign Zehpw6[0] = (~(Gbzhu6 & Nbzhu6));
assign Nbzhu6 = (~(T8yhu6 & Zazhu6));
assign T8yhu6 = (~(O9yhu6 | U5yhu6));
assign O9yhu6 = (Fnnhu6 & Ubzhu6);
assign Ubzhu6 = (Jayhu6 | Cayhu6);
assign Cayhu6 = (Bczhu6 & Ighpw6[4]);
assign Bczhu6 = (~(Ujyhu6 | Zwyhu6));
assign Gbzhu6 = (~(U5yhu6 & Iczhu6));
assign Iczhu6 = (~(Pczhu6 & Wczhu6));
assign Wczhu6 = (Ddzhu6 & Kdzhu6);
assign Kdzhu6 = (~(X9zhu6 | A1zhu6));
assign X9zhu6 = (Rdzhu6 & Iyyhu6);
assign Rdzhu6 = (~(Sbyhu6 | Ighpw6[0]));
assign Sbyhu6 = (Ydzhu6 & Fezhu6);
assign Fezhu6 = (Mdhpw6[1] & Mezhu6);
assign Mezhu6 = (Iahpw6[8] | Iahpw6[7]);
assign Ydzhu6 = (Tezhu6 & Pinhu6);
assign Ddzhu6 = (Afzhu6 & Iryhu6);
assign Iryhu6 = (~(Hfzhu6 & M7zhu6));
assign Hfzhu6 = (!T7zhu6);
assign T7zhu6 = (~(Ofzhu6 & Vfzhu6));
assign Vfzhu6 = (~(Cgzhu6 & Jgzhu6));
assign Jgzhu6 = (~(Ulnhu6 | Mdhpw6[1]));
assign Cgzhu6 = (~(Qgzhu6 | R7yhu6));
assign Afzhu6 = (~(Ziyhu6 & Ighpw6[4]));
assign Ziyhu6 = (~(Y7yhu6 | Zazhu6));
assign Pczhu6 = (Xgzhu6 & J9zhu6);
assign J9zhu6 = (Ehzhu6 & Lhzhu6);
assign Lhzhu6 = (~(Mdhpw6[3] & Agyhu6));
assign Ehzhu6 = (Shzhu6 & Ftyhu6);
assign Ftyhu6 = (~(Zhzhu6 & Ighpw6[2]));
assign Zhzhu6 = (~(Deyhu6 | Ighpw6[4]));
assign Shzhu6 = (~(Iyyhu6 & Gizhu6));
assign Gizhu6 = (~(Deyhu6 & Nizhu6));
assign Nizhu6 = (C9zhu6 | Mdhpw6[3]);
assign Xgzhu6 = (Uizhu6 & Bjzhu6);
assign Bjzhu6 = (~(Swyhu6 & Zazhu6));
assign Swyhu6 = (Ijzhu6 & Ighpw6[2]);
assign Uizhu6 = (~(Mdhpw6[3] & Pjzhu6));
assign Pjzhu6 = (~(Wjzhu6 & Dkzhu6));
assign Dkzhu6 = (~(Kkzhu6 | Hgyhu6));
assign Hgyhu6 = (Rkzhu6 & Zazhu6);
assign Kkzhu6 = (~(Tfyhu6 & Wryhu6));
assign Wryhu6 = (~(Ykzhu6 & Epyhu6));
assign Ykzhu6 = (~(Vuyhu6 | Deyhu6));
assign Tfyhu6 = (~(Rkzhu6 & Ighpw6[0]));
assign Rkzhu6 = (Flzhu6 & Epyhu6);
assign Flzhu6 = (~(Vuyhu6 | Ighpw6[1]));
assign Wjzhu6 = (Mlzhu6 & Tlzhu6);
assign Tlzhu6 = (~(M7zhu6 & Amzhu6));
assign M7zhu6 = (Hmzhu6 & Omzhu6);
assign Hmzhu6 = (~(Wdyhu6 | Vmzhu6));
assign Mlzhu6 = (Cnzhu6 & Joyhu6);
assign Cnzhu6 = (~(U4zhu6 & Jnzhu6));
assign Jnzhu6 = (~(Hknhu6 & Amzhu6));
assign Amzhu6 = (~(Mdhpw6[2] & Qnzhu6));
assign U4zhu6 = (!Pryhu6);
assign Pryhu6 = (~(Xnzhu6 & Eozhu6));
assign Eozhu6 = (~(Vmzhu6 | Ighpw6[1]));
assign Xnzhu6 = (~(Zazhu6 | Wdyhu6));
assign Zazhu6 = (!Ighpw6[0]);
assign Pkhpw6[1] = (~(Lozhu6 & Sozhu6));
assign Sozhu6 = (~(Zozhu6 & Gpzhu6));
assign Zozhu6 = (~(Npzhu6 & Upzhu6));
assign Upzhu6 = (~(Bqzhu6 & Iqzhu6));
assign Bqzhu6 = (~(Pqzhu6 | Wqzhu6));
assign Lozhu6 = (~(Drzhu6 & Krzhu6));
assign Pkhpw6[0] = (~(Rrzhu6 & Yrzhu6));
assign Yrzhu6 = (~(Krzhu6 & Fszhu6));
assign Rrzhu6 = (~(Mszhu6 | Tszhu6));
assign Mszhu6 = (Atzhu6 & Iqzhu6);
assign Atzhu6 = (~(Sqhpw6[0] | Sqhpw6[1]));
assign Vnfpw6[7] = (Ppfpw6[13] & Ivfhu6);
assign Vnfpw6[6] = (Ppfpw6[12] & Ivfhu6);
assign Vnfpw6[5] = (Ppfpw6[11] & Ivfhu6);
assign Vnfpw6[4] = (Ppfpw6[10] & Ivfhu6);
assign Vnfpw6[3] = (Ppfpw6[9] & Ivfhu6);
assign Vnfpw6[2] = (Ppfpw6[8] & Ivfhu6);
assign Vnfpw6[1] = (Ppfpw6[7] & Ivfhu6);
assign Vnfpw6[0] = (Ppfpw6[6] & Ivfhu6);
assign R0ghu6 = (~(Htzhu6 & Otzhu6));
assign Otzhu6 = (~(Vtzhu6 & Cuzhu6));
assign Htzhu6 = (Juzhu6 | Quzhu6);
assign Tgfpw6[9] = (~(Xuzhu6 | Evzhu6));
assign Tgfpw6[8] = (~(Xuzhu6 | Lvzhu6));
assign Tgfpw6[7] = (~(Xuzhu6 | Svzhu6));
assign Tgfpw6[6] = (~(Xuzhu6 | Zvzhu6));
assign Tgfpw6[5] = (~(Xuzhu6 | Gwzhu6));
assign Tgfpw6[4] = (~(Xuzhu6 | Nwzhu6));
assign Tgfpw6[3] = (~(Xuzhu6 | Uwzhu6));
assign Tgfpw6[31] = (~(Xuzhu6 | Bxzhu6));
assign Tgfpw6[30] = (~(Xuzhu6 | Ixzhu6));
assign Tgfpw6[2] = (~(Xuzhu6 | Pxzhu6));
assign Tgfpw6[29] = (~(Xuzhu6 | Wxzhu6));
assign Tgfpw6[28] = (~(Xuzhu6 | Dyzhu6));
assign Tgfpw6[27] = (~(Kyzhu6 | Xuzhu6));
assign Tgfpw6[26] = (~(Ryzhu6 | Xuzhu6));
assign Tgfpw6[25] = (~(Yyzhu6 | Xuzhu6));
assign Tgfpw6[24] = (~(Fzzhu6 | Xuzhu6));
assign Tgfpw6[23] = (~(Mzzhu6 | Xuzhu6));
assign Tgfpw6[22] = (~(Tzzhu6 | Xuzhu6));
assign Tgfpw6[21] = (~(A00iu6 | Xuzhu6));
assign Tgfpw6[20] = (~(H00iu6 | Xuzhu6));
assign Tgfpw6[1] = (~(Xuzhu6 | O00iu6));
assign Tgfpw6[19] = (~(V00iu6 | Xuzhu6));
assign Tgfpw6[18] = (~(C10iu6 | Xuzhu6));
assign Tgfpw6[17] = (~(J10iu6 | Xuzhu6));
assign Tgfpw6[16] = (~(Q10iu6 | Xuzhu6));
assign Tgfpw6[15] = (~(X10iu6 | Xuzhu6));
assign Tgfpw6[14] = (~(Xuzhu6 | E20iu6));
assign Tgfpw6[13] = (~(L20iu6 | Xuzhu6));
assign Tgfpw6[12] = (~(Xuzhu6 | S20iu6));
assign Tgfpw6[11] = (~(Xuzhu6 | Z20iu6));
assign Tgfpw6[10] = (~(Xuzhu6 | G30iu6));
assign Tgfpw6[0] = (~(Xuzhu6 | N30iu6));
assign Mifpw6[9] = (~(Xuzhu6 | U30iu6));
assign Mifpw6[8] = (~(Xuzhu6 | B40iu6));
assign Mifpw6[7] = (~(Xuzhu6 | I40iu6));
assign Mifpw6[6] = (~(Xuzhu6 | P40iu6));
assign Mifpw6[5] = (~(Xuzhu6 | W40iu6));
assign Mifpw6[4] = (~(Xuzhu6 | D50iu6));
assign Mifpw6[3] = (~(Xuzhu6 | K50iu6));
assign Mifpw6[31] = (~(Xuzhu6 | R50iu6));
assign Mifpw6[30] = (~(Xuzhu6 | Y50iu6));
assign Mifpw6[2] = (~(Xuzhu6 | F60iu6));
assign Mifpw6[29] = (~(Xuzhu6 | M60iu6));
assign Mifpw6[28] = (~(Xuzhu6 | T60iu6));
assign Mifpw6[27] = (~(Xuzhu6 | A70iu6));
assign Mifpw6[26] = (~(Xuzhu6 | H70iu6));
assign Mifpw6[25] = (~(Xuzhu6 | O70iu6));
assign Mifpw6[24] = (~(Xuzhu6 | V70iu6));
assign Mifpw6[23] = (~(Xuzhu6 | C80iu6));
assign Mifpw6[22] = (~(Xuzhu6 | J80iu6));
assign Mifpw6[21] = (~(Xuzhu6 | Q80iu6));
assign Mifpw6[20] = (~(Xuzhu6 | X80iu6));
assign Mifpw6[1] = (~(Xuzhu6 | E90iu6));
assign Mifpw6[19] = (~(Xuzhu6 | L90iu6));
assign Mifpw6[18] = (~(Xuzhu6 | S90iu6));
assign Mifpw6[17] = (~(Xuzhu6 | Z90iu6));
assign Mifpw6[16] = (~(Xuzhu6 | Ga0iu6));
assign Mifpw6[15] = (~(Xuzhu6 | Na0iu6));
assign Mifpw6[14] = (~(Xuzhu6 | Ua0iu6));
assign Mifpw6[13] = (~(Xuzhu6 | Bb0iu6));
assign Mifpw6[12] = (~(Xuzhu6 | Ib0iu6));
assign Mifpw6[11] = (~(Xuzhu6 | Pb0iu6));
assign Mifpw6[10] = (~(Xuzhu6 | Wb0iu6));
assign Mifpw6[0] = (~(Xuzhu6 | Dc0iu6));
assign Xuzhu6 = (Kc0iu6 & Rc0iu6);
assign Rc0iu6 = (~(Yc0iu6 & Fd0iu6));
assign Yc0iu6 = (C0ehu6 & Md0iu6);
assign Kc0iu6 = (Td0iu6 | Ae0iu6);
assign Idfpw6[9] = (He0iu6 & Oe0iu6);
assign Idfpw6[8] = (~(Ve0iu6 | Cf0iu6));
assign Idfpw6[7] = (~(Jf0iu6 | Cf0iu6));
assign Idfpw6[6] = (Qf0iu6 & Oe0iu6);
assign Idfpw6[5] = (~(Xf0iu6 | Cf0iu6));
assign Idfpw6[4] = (~(Eg0iu6 | Cf0iu6));
assign Idfpw6[3] = (~(Lg0iu6 | Cf0iu6));
assign Idfpw6[30] = (~(Sg0iu6 | Cf0iu6));
assign Idfpw6[2] = (Zg0iu6 & Gh0iu6);
assign Zg0iu6 = (Nh0iu6 & Oe0iu6);
assign Nh0iu6 = (~(Uh0iu6 & H6ghu6));
assign Uh0iu6 = (Bi0iu6 & Ii0iu6);
assign Idfpw6[29] = (~(Pi0iu6 | Cf0iu6));
assign Idfpw6[28] = (~(Wi0iu6 | Cf0iu6));
assign Idfpw6[27] = (Dj0iu6 & Oe0iu6);
assign Idfpw6[26] = (Kj0iu6 & Oe0iu6);
assign Idfpw6[25] = (Rj0iu6 & Oe0iu6);
assign Idfpw6[24] = (~(Yj0iu6 | Cf0iu6));
assign Idfpw6[23] = (~(Fk0iu6 | Cf0iu6));
assign Idfpw6[22] = (~(Mk0iu6 | Cf0iu6));
assign Idfpw6[21] = (~(Tk0iu6 | Cf0iu6));
assign Idfpw6[20] = (~(Al0iu6 | Cf0iu6));
assign Idfpw6[1] = (~(Hl0iu6 | Cf0iu6));
assign Idfpw6[19] = (~(Ol0iu6 | Cf0iu6));
assign Idfpw6[18] = (~(Vl0iu6 | Cf0iu6));
assign Idfpw6[17] = (~(Cm0iu6 | Cf0iu6));
assign Idfpw6[16] = (~(Jm0iu6 | Cf0iu6));
assign Idfpw6[15] = (~(Qm0iu6 | Cf0iu6));
assign Idfpw6[14] = (~(Xm0iu6 | Cf0iu6));
assign Idfpw6[13] = (~(En0iu6 | Cf0iu6));
assign Idfpw6[12] = (~(Ln0iu6 | Cf0iu6));
assign Idfpw6[11] = (~(Sn0iu6 | Cf0iu6));
assign Idfpw6[10] = (~(Zn0iu6 | Cf0iu6));
assign Cf0iu6 = (!Oe0iu6);
assign Idfpw6[0] = (Go0iu6 & Oe0iu6);
assign Dqfhu6 = (H6ghu6 & No0iu6);
assign No0iu6 = (~(Uo0iu6 & Bp0iu6));
assign Bp0iu6 = (Ip0iu6 & Pp0iu6);
assign Pp0iu6 = (~(Wp0iu6 & Dq0iu6));
assign Dq0iu6 = (~(Kq0iu6 & Rq0iu6));
assign Rq0iu6 = (~(Yq0iu6 & Fr0iu6));
assign Fr0iu6 = (~(Mr0iu6 | Tr0iu6));
assign Yq0iu6 = (~(As0iu6 | Hs0iu6));
assign Ip0iu6 = (~(C0ehu6 & Os0iu6));
assign Os0iu6 = (Vs0iu6 | Ct0iu6);
assign Ct0iu6 = (vis_apsr_o[1] & Jt0iu6);
assign Jt0iu6 = (~(Qt0iu6 & Xt0iu6));
assign Xt0iu6 = (Eu0iu6 | Cyfpw6[7]);
assign Qt0iu6 = (Mr0iu6 | Cyfpw6[3]);
assign Uo0iu6 = (Lu0iu6 & Su0iu6);
assign Su0iu6 = (Zu0iu6 | Cyfpw6[4]);
assign Eblhu6 = (Gv0iu6 & Rrlhu6);
assign Gv0iu6 = (Nv0iu6 ? Tzdpw6 : vis_pc_o[23]);
assign Lclhu6 = (Uv0iu6 & Kqlhu6);
assign Uv0iu6 = (Nv0iu6 ? A0epw6 : vis_pc_o[24]);
assign Sdlhu6 = (Bw0iu6 & Dplhu6);
assign Bw0iu6 = (Nv0iu6 ? H0epw6 : vis_pc_o[25]);
assign Zelhu6 = (Iw0iu6 & Wnlhu6);
assign Iw0iu6 = (Nv0iu6 ? O0epw6 : vis_pc_o[26]);
assign Gglhu6 = (Pw0iu6 & Pmlhu6);
assign Pw0iu6 = (Nv0iu6 ? V0epw6 : vis_pc_o[27]);
assign Nhlhu6 = (Ww0iu6 & Illhu6);
assign Ww0iu6 = (Nv0iu6 ? Dx0iu6 : vis_pc_o[28]);
assign Uilhu6 = (Kx0iu6 & Bklhu6);
assign Kx0iu6 = (Nv0iu6 ? Rx0iu6 : vis_pc_o[29]);
assign Knmhu6 = (Yx0iu6 | G4hpw6[0]);
assign Romhu6 = (Yx0iu6 | G4hpw6[1]);
assign Ypmhu6 = (Yx0iu6 | G4hpw6[2]);
assign Frmhu6 = (Yx0iu6 | G4hpw6[3]);
assign Gwhhu6 = (Fy0iu6 & A4khu6);
assign Fy0iu6 = (My0iu6 & Ty0iu6);
assign Oxhhu6 = (Az0iu6 & S2khu6);
assign Az0iu6 = (Ty0iu6 ? Hz0iu6 : vis_pc_o[0]);
assign Wyhhu6 = (Oz0iu6 & K1khu6);
assign Oz0iu6 = (Ty0iu6 ? Tugpw6[0] : vis_pc_o[1]);
assign E0ihu6 = (Vz0iu6 & C0khu6);
assign Vz0iu6 = (Ty0iu6 ? Tugpw6[1] : vis_pc_o[2]);
assign M1ihu6 = (C01iu6 & Uyjhu6);
assign C01iu6 = (Ty0iu6 ? Tugpw6[2] : vis_pc_o[3]);
assign U2ihu6 = (J01iu6 & Mxjhu6);
assign J01iu6 = (Ty0iu6 ? Tugpw6[3] : vis_pc_o[4]);
assign C4ihu6 = (Q01iu6 & Ewjhu6);
assign Q01iu6 = (Ty0iu6 ? Tugpw6[4] : vis_pc_o[5]);
assign K5ihu6 = (X01iu6 & Wujhu6);
assign X01iu6 = (Ty0iu6 ? Tugpw6[5] : vis_pc_o[6]);
assign S6ihu6 = (E11iu6 & Otjhu6);
assign E11iu6 = (Ty0iu6 ? Tugpw6[6] : vis_pc_o[7]);
assign Msmhu6 = (Yx0iu6 | G4hpw6[4]);
assign A8ihu6 = (L11iu6 & Gsjhu6);
assign L11iu6 = (Ty0iu6 ? Tugpw6[7] : vis_pc_o[8]);
assign I9ihu6 = (S11iu6 & Yqjhu6);
assign S11iu6 = (Ty0iu6 ? Tugpw6[8] : vis_pc_o[9]);
assign Qaihu6 = (Z11iu6 & Qpjhu6);
assign Z11iu6 = (Ty0iu6 ? Tugpw6[9] : vis_pc_o[10]);
assign Ybihu6 = (G21iu6 & Iojhu6);
assign G21iu6 = (Ty0iu6 ? Ixdpw6 : vis_pc_o[11]);
assign Gdihu6 = (N21iu6 & Anjhu6);
assign N21iu6 = (Ty0iu6 ? Tugpw6[11] : vis_pc_o[12]);
assign Oeihu6 = (U21iu6 & Sljhu6);
assign U21iu6 = (Ty0iu6 ? Tugpw6[12] : vis_pc_o[13]);
assign Wfihu6 = (B31iu6 & Kkjhu6);
assign B31iu6 = (Ty0iu6 ? Tugpw6[13] : vis_pc_o[14]);
assign Ehihu6 = (I31iu6 & Cjjhu6);
assign I31iu6 = (Ty0iu6 ? Pxdpw6 : vis_pc_o[15]);
assign Miihu6 = (P31iu6 & Uhjhu6);
assign P31iu6 = (Ty0iu6 ? Wxdpw6 : vis_pc_o[16]);
assign Ujihu6 = (W31iu6 & Mgjhu6);
assign W31iu6 = (Ty0iu6 ? Dydpw6 : vis_pc_o[17]);
assign Clihu6 = (D41iu6 & Efjhu6);
assign D41iu6 = (Ty0iu6 ? Kydpw6 : vis_pc_o[18]);
assign Kmihu6 = (K41iu6 & Wdjhu6);
assign K41iu6 = (Ty0iu6 ? Rydpw6 : vis_pc_o[19]);
assign Snihu6 = (R41iu6 & Ocjhu6);
assign R41iu6 = (Ty0iu6 ? Yydpw6 : vis_pc_o[20]);
assign Apihu6 = (Y41iu6 & Gbjhu6);
assign Y41iu6 = (Ty0iu6 ? Fzdpw6 : vis_pc_o[21]);
assign Iqihu6 = (F51iu6 & Y9jhu6);
assign F51iu6 = (Ty0iu6 ? Mzdpw6 : vis_pc_o[22]);
assign Qrihu6 = (M51iu6 & Q8jhu6);
assign M51iu6 = (Ty0iu6 ? Tzdpw6 : vis_pc_o[23]);
assign Ysihu6 = (T51iu6 & I7jhu6);
assign T51iu6 = (Ty0iu6 ? A0epw6 : vis_pc_o[24]);
assign Guihu6 = (A61iu6 & A6jhu6);
assign A61iu6 = (Ty0iu6 ? H0epw6 : vis_pc_o[25]);
assign Ovihu6 = (H61iu6 & S4jhu6);
assign H61iu6 = (Ty0iu6 ? O0epw6 : vis_pc_o[26]);
assign Wwihu6 = (O61iu6 & K3jhu6);
assign O61iu6 = (Ty0iu6 ? V0epw6 : vis_pc_o[27]);
assign Eyihu6 = (V61iu6 & C2jhu6);
assign V61iu6 = (Ty0iu6 ? Dx0iu6 : vis_pc_o[28]);
assign Mzihu6 = (C71iu6 & U0jhu6);
assign C71iu6 = (Ty0iu6 ? Rx0iu6 : vis_pc_o[29]);
assign Ttmhu6 = (V5hpw6[0] & J71iu6);
assign Avmhu6 = (V5hpw6[1] & Q71iu6);
assign Q71iu6 = (~(X71iu6 & Nv0iu6));
assign I5khu6 = (E81iu6 | Aygpw6[0]);
assign Q6khu6 = (E81iu6 | Aygpw6[1]);
assign Y7khu6 = (E81iu6 | Aygpw6[2]);
assign G9khu6 = (E81iu6 | Aygpw6[3]);
assign Oakhu6 = (E81iu6 | Aygpw6[4]);
assign Wbkhu6 = (Pzgpw6[0] & J71iu6);
assign Edkhu6 = (Pzgpw6[1] & L81iu6);
assign L81iu6 = (~(X71iu6 & Ty0iu6));
assign Ufkhu6 = (S81iu6 & Dmmhu6);
assign S81iu6 = (My0iu6 & Nv0iu6);
assign Chkhu6 = (Z81iu6 & Wkmhu6);
assign Z81iu6 = (Nv0iu6 ? Hz0iu6 : vis_pc_o[0]);
assign Kikhu6 = (G91iu6 & Pjmhu6);
assign G91iu6 = (Nv0iu6 ? Tugpw6[0] : vis_pc_o[1]);
assign Sjkhu6 = (N91iu6 & Iimhu6);
assign N91iu6 = (Nv0iu6 ? Tugpw6[1] : vis_pc_o[2]);
assign Alkhu6 = (U91iu6 & Bhmhu6);
assign U91iu6 = (Nv0iu6 ? Tugpw6[2] : vis_pc_o[3]);
assign Imkhu6 = (Ba1iu6 & Ufmhu6);
assign Ba1iu6 = (Nv0iu6 ? Tugpw6[3] : vis_pc_o[4]);
assign Qnkhu6 = (Ia1iu6 & Nemhu6);
assign Ia1iu6 = (Nv0iu6 ? Tugpw6[4] : vis_pc_o[5]);
assign Yokhu6 = (Pa1iu6 & Gdmhu6);
assign Pa1iu6 = (Nv0iu6 ? Tugpw6[5] : vis_pc_o[6]);
assign Gqkhu6 = (Wa1iu6 & Zbmhu6);
assign Wa1iu6 = (Nv0iu6 ? Tugpw6[6] : vis_pc_o[7]);
assign Orkhu6 = (Db1iu6 & Samhu6);
assign Db1iu6 = (Nv0iu6 ? Tugpw6[7] : vis_pc_o[8]);
assign Wskhu6 = (Kb1iu6 & L9mhu6);
assign Kb1iu6 = (Nv0iu6 ? Tugpw6[8] : vis_pc_o[9]);
assign Eukhu6 = (Rb1iu6 & E8mhu6);
assign Rb1iu6 = (Nv0iu6 ? Tugpw6[9] : vis_pc_o[10]);
assign Mvkhu6 = (Yb1iu6 & X6mhu6);
assign Yb1iu6 = (Nv0iu6 ? Ixdpw6 : vis_pc_o[11]);
assign Uwkhu6 = (Fc1iu6 & Q5mhu6);
assign Fc1iu6 = (Nv0iu6 ? Tugpw6[11] : vis_pc_o[12]);
assign Cykhu6 = (Mc1iu6 & J4mhu6);
assign Mc1iu6 = (Nv0iu6 ? Tugpw6[12] : vis_pc_o[13]);
assign Kzkhu6 = (Tc1iu6 & C3mhu6);
assign Tc1iu6 = (Nv0iu6 ? Tugpw6[13] : vis_pc_o[14]);
assign S0lhu6 = (Ad1iu6 & V1mhu6);
assign Ad1iu6 = (Nv0iu6 ? Pxdpw6 : vis_pc_o[15]);
assign A2lhu6 = (Hd1iu6 & O0mhu6);
assign Hd1iu6 = (Nv0iu6 ? Wxdpw6 : vis_pc_o[16]);
assign I3lhu6 = (Od1iu6 & Hzlhu6);
assign Od1iu6 = (Nv0iu6 ? Dydpw6 : vis_pc_o[17]);
assign Q4lhu6 = (Vd1iu6 & Aylhu6);
assign Vd1iu6 = (Nv0iu6 ? Kydpw6 : vis_pc_o[18]);
assign Y5lhu6 = (Ce1iu6 & Twlhu6);
assign Ce1iu6 = (Nv0iu6 ? Rydpw6 : vis_pc_o[19]);
assign G7lhu6 = (Je1iu6 & Mvlhu6);
assign Je1iu6 = (Nv0iu6 ? Yydpw6 : vis_pc_o[20]);
assign O8lhu6 = (Qe1iu6 & Fulhu6);
assign Qe1iu6 = (Nv0iu6 ? Fzdpw6 : vis_pc_o[21]);
assign W9lhu6 = (Xe1iu6 & Yslhu6);
assign Xe1iu6 = (Nv0iu6 ? Mzdpw6 : vis_pc_o[22]);
assign R9ohu6 = (Ty0iu6 ? Ef1iu6 : vis_pc_o[30]);
assign M9ohu6 = (Nv0iu6 ? Ef1iu6 : vis_pc_o[30]);
assign X3yhu6 = (Sf1iu6 ? X0ohu6 : Lf1iu6);
assign Q3yhu6 = (~(Zf1iu6 & Gg1iu6));
assign Gg1iu6 = (Ng1iu6 | Ug1iu6);
assign Ug1iu6 = (!Bh1iu6);
assign Zf1iu6 = (~(Ih1iu6 | Ph1iu6));
assign Ih1iu6 = (Fanhu6 & Wh1iu6);
assign Wh1iu6 = (~(Iahpw6[1] & Di1iu6));
assign J3yhu6 = (~(Ki1iu6 & Ri1iu6));
assign Ri1iu6 = (~(Yi1iu6 & Fj1iu6));
assign Yi1iu6 = (~(Ofzhu6 | Mdhpw6[0]));
assign Ki1iu6 = (~(Jdnhu6 & Mj1iu6));
assign Mj1iu6 = (~(Iahpw6[2] & Di1iu6));
assign C3yhu6 = (~(Tj1iu6 & Ak1iu6));
assign Ak1iu6 = (Hk1iu6 & Ok1iu6);
assign Ok1iu6 = (~(Uthpw6[7] & Vk1iu6));
assign Hk1iu6 = (~(Cl1iu6 & Jdnhu6));
assign Tj1iu6 = (Jl1iu6 & Ql1iu6);
assign Ql1iu6 = (~(Iahpw6[6] & Xl1iu6));
assign Jl1iu6 = (~(Iahpw6[7] & Z4yhu6));
assign V2yhu6 = (Em1iu6 ? Iahpw6[30] : Shhpw6[31]);
assign O2yhu6 = (Sm1iu6 ? Lm1iu6 : Jshpw6[31]);
assign H2yhu6 = (~(Zm1iu6 & Gn1iu6));
assign Gn1iu6 = (Nn1iu6 & Un1iu6);
assign Un1iu6 = (~(Bo1iu6 & Jshpw6[31]));
assign Nn1iu6 = (Io1iu6 & Po1iu6);
assign Io1iu6 = (~(Wo1iu6 & Dp1iu6));
assign Dp1iu6 = (~(Kp1iu6 & Rp1iu6));
assign Rp1iu6 = (Yp1iu6 & Fq1iu6);
assign Fq1iu6 = (Mq1iu6 & Tq1iu6);
assign Tq1iu6 = (~(Ar1iu6 & Fkfpw6[31]));
assign Mq1iu6 = (Hr1iu6 & Or1iu6);
assign Or1iu6 = (~(Ligpw6[28] & Vr1iu6));
assign Hr1iu6 = (~(Engpw6[28] & Cs1iu6));
assign Yp1iu6 = (Js1iu6 & Qs1iu6);
assign Qs1iu6 = (~(Akgpw6[28] & Xs1iu6));
assign Js1iu6 = (Et1iu6 & Lt1iu6);
assign Lt1iu6 = (~(HRDATA[31] & St1iu6));
assign Et1iu6 = (~(E1hpw6[31] & Zt1iu6));
assign Kp1iu6 = (Gu1iu6 & Nu1iu6);
assign Nu1iu6 = (Uu1iu6 & Bv1iu6);
assign Bv1iu6 = (~(Iv1iu6 & vis_pc_o[30]));
assign Uu1iu6 = (Pv1iu6 & Wv1iu6);
assign Wv1iu6 = (~(Plgpw6[28] & Dw1iu6));
assign Pv1iu6 = (~(K7hpw6[31] & Kw1iu6));
assign Gu1iu6 = (Rw1iu6 & Yw1iu6);
assign Zm1iu6 = (Fx1iu6 & Mx1iu6);
assign Mx1iu6 = (~(ECOREVNUM[23] & Tx1iu6));
assign Fx1iu6 = (~(Uthpw6[31] & Sf1iu6));
assign A2yhu6 = (~(Ay1iu6 & Hy1iu6));
assign Hy1iu6 = (Oy1iu6 & Vy1iu6);
assign Oy1iu6 = (Cz1iu6 & Jz1iu6);
assign Jz1iu6 = (~(Uthpw6[31] & Vk1iu6));
assign Cz1iu6 = (~(ECOREVNUM[27] & Qz1iu6));
assign Ay1iu6 = (Xz1iu6 & E02iu6);
assign E02iu6 = (~(Iahpw6[30] & Xl1iu6));
assign Xz1iu6 = (L02iu6 | Jayhu6);
assign Jayhu6 = (!Mdhpw6[3]);
assign T1yhu6 = (~(S02iu6 & Z02iu6));
assign Z02iu6 = (G12iu6 & Vy1iu6);
assign Vy1iu6 = (~(Zbhpw6[30] & Cl1iu6));
assign G12iu6 = (N12iu6 & U12iu6);
assign U12iu6 = (~(Uthpw6[30] & Vk1iu6));
assign N12iu6 = (~(ECOREVNUM[26] & Qz1iu6));
assign S02iu6 = (B22iu6 & I22iu6);
assign I22iu6 = (~(Iahpw6[29] & Xl1iu6));
assign B22iu6 = (~(Iahpw6[30] & Z4yhu6));
assign M1yhu6 = (~(P22iu6 & W22iu6));
assign W22iu6 = (D32iu6 & K32iu6);
assign K32iu6 = (~(ECOREVNUM[25] & Qz1iu6));
assign D32iu6 = (R32iu6 & Y32iu6);
assign Y32iu6 = (~(F42iu6 & Cl1iu6));
assign F42iu6 = (Gwnhu6 & M42iu6);
assign M42iu6 = (~(Zbhpw6[28] & T42iu6));
assign T42iu6 = (A52iu6 | W9ohu6);
assign R32iu6 = (~(Uthpw6[29] & Vk1iu6));
assign P22iu6 = (H52iu6 & O52iu6);
assign O52iu6 = (~(Iahpw6[28] & Xl1iu6));
assign H52iu6 = (~(Iahpw6[29] & Z4yhu6));
assign F1yhu6 = (~(V52iu6 & C62iu6));
assign C62iu6 = (J62iu6 & Q62iu6);
assign Q62iu6 = (~(Cl1iu6 & Zbhpw6[28]));
assign J62iu6 = (X62iu6 & E72iu6);
assign E72iu6 = (~(Uthpw6[28] & Vk1iu6));
assign X62iu6 = (~(ECOREVNUM[24] & Qz1iu6));
assign Qz1iu6 = (!L72iu6);
assign V52iu6 = (S72iu6 & Z72iu6);
assign Z72iu6 = (~(Iahpw6[27] & Xl1iu6));
assign S72iu6 = (~(Iahpw6[28] & Z4yhu6));
assign Y0yhu6 = (~(G82iu6 & N82iu6));
assign N82iu6 = (U82iu6 & L72iu6);
assign U82iu6 = (~(Uthpw6[27] & Vk1iu6));
assign G82iu6 = (B92iu6 & I92iu6);
assign I92iu6 = (~(Iahpw6[26] & Xl1iu6));
assign B92iu6 = (~(Iahpw6[27] & Z4yhu6));
assign R0yhu6 = (~(P92iu6 & W92iu6));
assign W92iu6 = (Da2iu6 & Ka2iu6);
assign Ka2iu6 = (~(Uthpw6[26] & Vk1iu6));
assign Da2iu6 = (~(Zbhpw6[26] & Cl1iu6));
assign P92iu6 = (Ra2iu6 & Ya2iu6);
assign Ya2iu6 = (~(Iahpw6[25] & Xl1iu6));
assign Ra2iu6 = (~(Iahpw6[26] & Z4yhu6));
assign K0yhu6 = (~(Fb2iu6 & Mb2iu6));
assign Mb2iu6 = (Tb2iu6 & L72iu6);
assign Tb2iu6 = (~(Uthpw6[25] & Vk1iu6));
assign Fb2iu6 = (Ac2iu6 & Hc2iu6);
assign Hc2iu6 = (~(Iahpw6[24] & Xl1iu6));
assign Ac2iu6 = (~(Iahpw6[25] & Z4yhu6));
assign D0yhu6 = (~(Oc2iu6 & Vc2iu6));
assign Vc2iu6 = (Cd2iu6 & L72iu6);
assign Cd2iu6 = (~(Uthpw6[24] & Vk1iu6));
assign Oc2iu6 = (Jd2iu6 & Qd2iu6);
assign Qd2iu6 = (~(Iahpw6[23] & Xl1iu6));
assign Jd2iu6 = (~(Iahpw6[24] & Z4yhu6));
assign Wzxhu6 = (~(Xd2iu6 & Ee2iu6));
assign Ee2iu6 = (Le2iu6 & L72iu6);
assign Le2iu6 = (~(Uthpw6[23] & Vk1iu6));
assign Xd2iu6 = (Se2iu6 & Ze2iu6);
assign Ze2iu6 = (~(Iahpw6[22] & Xl1iu6));
assign Se2iu6 = (~(Iahpw6[23] & Z4yhu6));
assign Pzxhu6 = (~(Gf2iu6 & Nf2iu6));
assign Nf2iu6 = (~(Iahpw6[22] & Z4yhu6));
assign Gf2iu6 = (Uf2iu6 & Bg2iu6);
assign Bg2iu6 = (~(Uthpw6[22] & Vk1iu6));
assign Uf2iu6 = (~(Iahpw6[21] & Xl1iu6));
assign Izxhu6 = (~(Ig2iu6 & Pg2iu6));
assign Pg2iu6 = (Wg2iu6 & L72iu6);
assign Wg2iu6 = (~(Uthpw6[21] & Vk1iu6));
assign Ig2iu6 = (Dh2iu6 & Kh2iu6);
assign Kh2iu6 = (~(Iahpw6[20] & Xl1iu6));
assign Dh2iu6 = (~(Iahpw6[21] & Z4yhu6));
assign Bzxhu6 = (~(Rh2iu6 & Yh2iu6));
assign Yh2iu6 = (Fi2iu6 & L72iu6);
assign Fi2iu6 = (~(Uthpw6[20] & Vk1iu6));
assign Rh2iu6 = (Mi2iu6 & Ti2iu6);
assign Ti2iu6 = (~(Iahpw6[19] & Xl1iu6));
assign Mi2iu6 = (~(Iahpw6[20] & Z4yhu6));
assign Uyxhu6 = (~(Aj2iu6 & Hj2iu6));
assign Hj2iu6 = (~(Iahpw6[19] & Z4yhu6));
assign Aj2iu6 = (Oj2iu6 & Vj2iu6);
assign Vj2iu6 = (~(Uthpw6[19] & Vk1iu6));
assign Oj2iu6 = (~(Iahpw6[18] & Xl1iu6));
assign Nyxhu6 = (~(Ck2iu6 & Jk2iu6));
assign Jk2iu6 = (~(Iahpw6[18] & Z4yhu6));
assign Ck2iu6 = (Qk2iu6 & Xk2iu6);
assign Xk2iu6 = (~(Uthpw6[18] & Vk1iu6));
assign Qk2iu6 = (~(Iahpw6[17] & Xl1iu6));
assign Gyxhu6 = (~(El2iu6 & Ll2iu6));
assign Ll2iu6 = (~(Iahpw6[17] & Z4yhu6));
assign El2iu6 = (Sl2iu6 & Zl2iu6);
assign Zl2iu6 = (~(Uthpw6[17] & Vk1iu6));
assign Sl2iu6 = (~(Iahpw6[16] & Xl1iu6));
assign Zxxhu6 = (~(Gm2iu6 & Nm2iu6));
assign Nm2iu6 = (Um2iu6 & L72iu6);
assign Um2iu6 = (~(Uthpw6[16] & Vk1iu6));
assign Gm2iu6 = (Bn2iu6 & In2iu6);
assign In2iu6 = (~(Iahpw6[15] & Xl1iu6));
assign Bn2iu6 = (~(Iahpw6[16] & Z4yhu6));
assign Sxxhu6 = (~(Pn2iu6 & Wn2iu6));
assign Wn2iu6 = (~(Iahpw6[15] & Z4yhu6));
assign Pn2iu6 = (Do2iu6 & Ko2iu6);
assign Ko2iu6 = (~(Uthpw6[15] & Vk1iu6));
assign Do2iu6 = (~(Iahpw6[14] & Xl1iu6));
assign Lxxhu6 = (~(Ro2iu6 & Yo2iu6));
assign Yo2iu6 = (~(Iahpw6[14] & Z4yhu6));
assign Ro2iu6 = (Fp2iu6 & Mp2iu6);
assign Mp2iu6 = (~(Uthpw6[14] & Vk1iu6));
assign Fp2iu6 = (~(Iahpw6[13] & Xl1iu6));
assign Exxhu6 = (~(Tp2iu6 & Aq2iu6));
assign Aq2iu6 = (~(Iahpw6[13] & Z4yhu6));
assign Tp2iu6 = (Hq2iu6 & Oq2iu6);
assign Oq2iu6 = (~(Uthpw6[13] & Vk1iu6));
assign Hq2iu6 = (~(Iahpw6[12] & Xl1iu6));
assign Xwxhu6 = (~(Vq2iu6 & Cr2iu6));
assign Cr2iu6 = (Jr2iu6 & L72iu6);
assign Jr2iu6 = (~(Uthpw6[12] & Vk1iu6));
assign Vq2iu6 = (Qr2iu6 & Xr2iu6);
assign Xr2iu6 = (~(Iahpw6[11] & Xl1iu6));
assign Qr2iu6 = (~(Iahpw6[12] & Z4yhu6));
assign Qwxhu6 = (~(Es2iu6 & Ls2iu6));
assign Ls2iu6 = (~(Iahpw6[11] & Z4yhu6));
assign Es2iu6 = (Ss2iu6 & Zs2iu6);
assign Zs2iu6 = (~(Uthpw6[11] & Vk1iu6));
assign Ss2iu6 = (~(Iahpw6[10] & Xl1iu6));
assign Jwxhu6 = (~(Gt2iu6 & Nt2iu6));
assign Nt2iu6 = (Ut2iu6 & L72iu6);
assign Ut2iu6 = (~(Uthpw6[10] & Vk1iu6));
assign Gt2iu6 = (Bu2iu6 & Iu2iu6);
assign Iu2iu6 = (~(Iahpw6[9] & Xl1iu6));
assign Bu2iu6 = (~(Iahpw6[10] & Z4yhu6));
assign Cwxhu6 = (~(Pu2iu6 & Wu2iu6));
assign Wu2iu6 = (~(Iahpw6[9] & Z4yhu6));
assign Pu2iu6 = (Dv2iu6 & Kv2iu6);
assign Kv2iu6 = (~(Uthpw6[9] & Vk1iu6));
assign Dv2iu6 = (~(Iahpw6[8] & Xl1iu6));
assign Vvxhu6 = (~(Rv2iu6 & Yv2iu6));
assign Yv2iu6 = (~(Iahpw6[8] & Z4yhu6));
assign Rv2iu6 = (Fw2iu6 & Mw2iu6);
assign Mw2iu6 = (~(Uthpw6[8] & Vk1iu6));
assign Fw2iu6 = (~(Iahpw6[7] & Xl1iu6));
assign Ovxhu6 = (Tw2iu6 ? Mdhpw6[3] : SWDITMS);
assign Tw2iu6 = (Ax2iu6 & Hx2iu6);
assign Hx2iu6 = (Ox2iu6 & Vx2iu6);
assign Ox2iu6 = (~(Cy2iu6 & Ujyhu6));
assign Cy2iu6 = (Jy2iu6 | Qy2iu6);
assign Qy2iu6 = (Ighpw6[1] ? Iyyhu6 : Xy2iu6);
assign Xy2iu6 = (Ez2iu6 & Lz2iu6);
assign Lz2iu6 = (~(Wdyhu6 & Sz2iu6));
assign Sz2iu6 = (Mdhpw6[0] | Ighpw6[0]);
assign Jy2iu6 = (~(Zz2iu6 & G03iu6));
assign G03iu6 = (~(N03iu6 & Ighpw6[2]));
assign N03iu6 = (Gjyhu6 & Eiyhu6);
assign Zz2iu6 = (Deyhu6 | Ighpw6[3]);
assign Ax2iu6 = (U03iu6 & B13iu6);
assign B13iu6 = (L02iu6 | Mdhpw6[0]);
assign Hvxhu6 = (W13iu6 ? P13iu6 : I13iu6);
assign I13iu6 = (D23iu6 & K23iu6);
assign K23iu6 = (R23iu6 & Y23iu6);
assign Y23iu6 = (~(Iahpw6[29] | Iahpw6[30]));
assign R23iu6 = (~(Iahpw6[27] | Iahpw6[28]));
assign D23iu6 = (F33iu6 & M33iu6);
assign M33iu6 = (~(Iahpw6[25] | Iahpw6[26]));
assign F33iu6 = (~(Iahpw6[23] | Iahpw6[24]));
assign Avxhu6 = (W13iu6 ? A43iu6 : T33iu6);
assign A43iu6 = (!Omdpw6);
assign Tuxhu6 = (Em1iu6 ? H43iu6 : Cjhpw6[3]);
assign H43iu6 = (~(Omdpw6 & O43iu6));
assign Muxhu6 = (V43iu6 ? Lznhu6 : Dtnhu6);
assign V43iu6 = (~(Npzhu6 | Gpzhu6));
assign Fuxhu6 = (~(C53iu6 ^ G2ohu6));
assign Ytxhu6 = (Q53iu6 ? Punhu6 : J53iu6);
assign Q53iu6 = (~(Rrnhu6 | G2ohu6));
assign J53iu6 = (!W9ohu6);
assign Rtxhu6 = (~(X53iu6 & E63iu6));
assign E63iu6 = (~(Rgnhu6 & L63iu6));
assign L63iu6 = (~(S63iu6 & Fmyhu6));
assign S63iu6 = (~(Z63iu6 | G73iu6));
assign G73iu6 = (~(N73iu6 | R7yhu6));
assign Ktxhu6 = (U73iu6 ? Mmyhu6 : Ubnhu6);
assign U73iu6 = (B83iu6 & Mdhpw6[0]);
assign B83iu6 = (~(N5yhu6 | I83iu6));
assign Dtxhu6 = (~(P83iu6 & W83iu6));
assign W83iu6 = (D93iu6 & K93iu6);
assign K93iu6 = (~(Uthpw6[6] & Vk1iu6));
assign D93iu6 = (R93iu6 & L72iu6);
assign R93iu6 = (~(Y93iu6 & Pinhu6));
assign P83iu6 = (Fa3iu6 & Ma3iu6);
assign Ma3iu6 = (~(Iahpw6[6] & Z4yhu6));
assign Fa3iu6 = (Ta3iu6 & Ab3iu6);
assign Ab3iu6 = (~(Ubnhu6 & Cl1iu6));
assign Ta3iu6 = (~(Iahpw6[5] & Xl1iu6));
assign Wsxhu6 = (~(Hb3iu6 & Ob3iu6));
assign Ob3iu6 = (Vb3iu6 & Cc3iu6);
assign Cc3iu6 = (~(Cl1iu6 & Fanhu6));
assign Vb3iu6 = (Jc3iu6 & L72iu6);
assign Jc3iu6 = (~(Uthpw6[5] & Vk1iu6));
assign Hb3iu6 = (Qc3iu6 & Xc3iu6);
assign Xc3iu6 = (~(Iahpw6[4] & Xl1iu6));
assign Qc3iu6 = (~(Iahpw6[5] & Z4yhu6));
assign Psxhu6 = (~(Ed3iu6 & Ld3iu6));
assign Ld3iu6 = (Sd3iu6 & L72iu6);
assign Sd3iu6 = (~(Uthpw6[4] & Vk1iu6));
assign Ed3iu6 = (Zd3iu6 & Ge3iu6);
assign Ge3iu6 = (~(Iahpw6[3] & Xl1iu6));
assign Zd3iu6 = (~(Iahpw6[4] & Z4yhu6));
assign Isxhu6 = (W13iu6 ? N3nhu6 : Ne3iu6);
assign Ne3iu6 = (Iahpw6[3] & Ue3iu6);
assign Ue3iu6 = (~(T33iu6 & Bf3iu6));
assign Bf3iu6 = (~(If3iu6 & Iahpw6[4]));
assign If3iu6 = (Iahpw6[5] & Iahpw6[6]);
assign T33iu6 = (Pf3iu6 | Iahpw6[4]);
assign Pf3iu6 = (Iahpw6[5] | Iahpw6[6]);
assign Bsxhu6 = (~(Wf3iu6 & Dg3iu6));
assign Dg3iu6 = (~(Iahpw6[3] & Z4yhu6));
assign Wf3iu6 = (Kg3iu6 & Rg3iu6);
assign Rg3iu6 = (~(Uthpw6[3] & Vk1iu6));
assign Kg3iu6 = (~(Xl1iu6 & Iahpw6[2]));
assign Urxhu6 = (~(Yg3iu6 & Fh3iu6));
assign Fh3iu6 = (Mh3iu6 & L72iu6);
assign Mh3iu6 = (~(Uthpw6[2] & Vk1iu6));
assign Yg3iu6 = (Th3iu6 & Ai3iu6);
assign Ai3iu6 = (~(Xl1iu6 & Iahpw6[1]));
assign Th3iu6 = (~(Iahpw6[2] & Z4yhu6));
assign Nrxhu6 = (~(Hi3iu6 & Oi3iu6));
assign Oi3iu6 = (~(Vi3iu6 & B7nhu6));
assign Vi3iu6 = (Cj3iu6 & L02iu6);
assign Cj3iu6 = (~(Vx2iu6 & Jj3iu6));
assign Jj3iu6 = (~(A1zhu6 & Qj3iu6));
assign Qj3iu6 = (Hknhu6 | K7yhu6);
assign K7yhu6 = (!Xj3iu6);
assign Hi3iu6 = (~(Q8nhu6 & Ek3iu6));
assign Ek3iu6 = (~(Iahpw6[3] & Di1iu6));
assign Grxhu6 = (~(Lk3iu6 & Sk3iu6));
assign Sk3iu6 = (Zk3iu6 & Gl3iu6);
assign Gl3iu6 = (~(Q8nhu6 & Cl1iu6));
assign Zk3iu6 = (Nl3iu6 & L72iu6);
assign Nl3iu6 = (~(Uthpw6[1] & Vk1iu6));
assign Lk3iu6 = (Ul3iu6 & Bm3iu6);
assign Bm3iu6 = (~(Iahpw6[0] & Xl1iu6));
assign Ul3iu6 = (~(Iahpw6[1] & Z4yhu6));
assign Zqxhu6 = (~(Im3iu6 & Pm3iu6));
assign Pm3iu6 = (Wm3iu6 & Dn3iu6);
assign Dn3iu6 = (~(B7nhu6 & Cl1iu6));
assign Cl1iu6 = (Kn3iu6 & Y93iu6);
assign Wm3iu6 = (Rn3iu6 & L72iu6);
assign L72iu6 = (~(Y93iu6 & O8zhu6));
assign Y93iu6 = (Yn3iu6 & Fmyhu6);
assign Rn3iu6 = (~(Uthpw6[0] & Vk1iu6));
assign Vk1iu6 = (Fo3iu6 & Mo3iu6);
assign Fo3iu6 = (~(I83iu6 | Yenhu6));
assign I83iu6 = (!N73iu6);
assign Im3iu6 = (To3iu6 & Ap3iu6);
assign Ap3iu6 = (~(Tonhu6 & Xl1iu6));
assign Xl1iu6 = (~(Z4yhu6 | Fmyhu6));
assign To3iu6 = (~(Iahpw6[0] & Z4yhu6));
assign Sqxhu6 = (W13iu6 ? Pinhu6 : Tonhu6);
assign W13iu6 = (~(Hp3iu6 & Op3iu6));
assign Op3iu6 = (~(Vp3iu6 | Mdhpw6[1]));
assign Hp3iu6 = (Mdhpw6[2] & Cq3iu6);
assign Lqxhu6 = (Jq3iu6 ? Zbhpw6[30] : Iahpw6[29]);
assign Eqxhu6 = (Em1iu6 ? Mdhpw6[2] : Cjhpw6[1]);
assign Xpxhu6 = (Em1iu6 ? Qq3iu6 : Cjhpw6[2]);
assign Qq3iu6 = (N3nhu6 & O43iu6);
assign Qpxhu6 = (Em1iu6 ? Mdhpw6[1] : Cjhpw6[0]);
assign Jpxhu6 = (Em1iu6 ? Iahpw6[0] : Shhpw6[1]);
assign Cpxhu6 = (Em1iu6 ? Iahpw6[1] : Shhpw6[2]);
assign Voxhu6 = (Em1iu6 ? Iahpw6[2] : Shhpw6[3]);
assign Ooxhu6 = (Em1iu6 ? Iahpw6[3] : Shhpw6[4]);
assign Hoxhu6 = (Em1iu6 ? Iahpw6[4] : Shhpw6[5]);
assign Aoxhu6 = (Em1iu6 ? Iahpw6[5] : Shhpw6[6]);
assign Tnxhu6 = (Em1iu6 ? Iahpw6[6] : Shhpw6[7]);
assign Mnxhu6 = (Em1iu6 ? Iahpw6[7] : Shhpw6[8]);
assign Fnxhu6 = (Em1iu6 ? Iahpw6[8] : Shhpw6[9]);
assign Ymxhu6 = (Em1iu6 ? Iahpw6[9] : Shhpw6[10]);
assign Rmxhu6 = (Em1iu6 ? Iahpw6[10] : Shhpw6[11]);
assign Kmxhu6 = (Em1iu6 ? Iahpw6[11] : Shhpw6[12]);
assign Dmxhu6 = (Em1iu6 ? Iahpw6[12] : Shhpw6[13]);
assign Wlxhu6 = (Em1iu6 ? Iahpw6[13] : Shhpw6[14]);
assign Plxhu6 = (Em1iu6 ? Iahpw6[14] : Shhpw6[15]);
assign Ilxhu6 = (Em1iu6 ? Iahpw6[15] : Shhpw6[16]);
assign Blxhu6 = (Em1iu6 ? Iahpw6[16] : Shhpw6[17]);
assign Ukxhu6 = (Em1iu6 ? Iahpw6[17] : Shhpw6[18]);
assign Nkxhu6 = (Em1iu6 ? Iahpw6[18] : Shhpw6[19]);
assign Gkxhu6 = (Em1iu6 ? Iahpw6[19] : Shhpw6[20]);
assign Zjxhu6 = (Em1iu6 ? Iahpw6[20] : Shhpw6[21]);
assign Sjxhu6 = (Em1iu6 ? Iahpw6[21] : Shhpw6[22]);
assign Ljxhu6 = (Em1iu6 ? Iahpw6[22] : Shhpw6[23]);
assign Ejxhu6 = (Em1iu6 ? Iahpw6[23] : Shhpw6[24]);
assign Xixhu6 = (Em1iu6 ? Iahpw6[24] : Shhpw6[25]);
assign Qixhu6 = (Em1iu6 ? Iahpw6[25] : Shhpw6[26]);
assign Jixhu6 = (Em1iu6 ? Iahpw6[26] : Shhpw6[27]);
assign Cixhu6 = (Em1iu6 ? Iahpw6[27] : Shhpw6[28]);
assign Vhxhu6 = (Em1iu6 ? Iahpw6[28] : Shhpw6[29]);
assign Ohxhu6 = (Em1iu6 ? Iahpw6[29] : Shhpw6[30]);
assign Hhxhu6 = (Em1iu6 ? Tonhu6 : Shhpw6[0]);
assign Ahxhu6 = (Em1iu6 ? Mdhpw6[0] : Iqnhu6);
assign Em1iu6 = (!C53iu6);
assign C53iu6 = (X53iu6 & O43iu6);
assign O43iu6 = (~(Xq3iu6 & G2ohu6));
assign Xq3iu6 = (Rrnhu6 & A52iu6);
assign X53iu6 = (Bh1iu6 | Ng1iu6);
assign Ng1iu6 = (~(Er3iu6 & Lr3iu6));
assign Lr3iu6 = (Sr3iu6 & P13iu6);
assign Sr3iu6 = (Ofzhu6 | Mdhpw6[0]);
assign Ofzhu6 = (!Vp3iu6);
assign Er3iu6 = (Ulnhu6 & Fj1iu6);
assign Bh1iu6 = (~(Zr3iu6 & Gs3iu6));
assign Gs3iu6 = (~(A52iu6 | W9ohu6));
assign Zr3iu6 = (Zbhpw6[28] & Gwnhu6);
assign Tgxhu6 = (Jq3iu6 ? B7nhu6 : Tonhu6);
assign Mgxhu6 = (Jq3iu6 ? Zbhpw6[26] : Iahpw6[25]);
assign Fgxhu6 = (Jq3iu6 ? Zbhpw6[28] : Iahpw6[27]);
assign Jq3iu6 = (~(Kn3iu6 & Tezhu6));
assign Kn3iu6 = (~(O8zhu6 | Pinhu6));
assign Yfxhu6 = (~(Ns3iu6 & Us3iu6));
assign Us3iu6 = (~(Zbhpw6[28] & Bt3iu6));
assign Bt3iu6 = (~(Gwnhu6 & A52iu6));
assign Ns3iu6 = (A52iu6 | Gwnhu6);
assign A52iu6 = (!Punhu6);
assign Rfxhu6 = (~(It3iu6 & Pt3iu6));
assign Pt3iu6 = (~(U5yhu6 & Wt3iu6));
assign Wt3iu6 = (Du3iu6 | Ku3iu6);
assign Ku3iu6 = (Mmyhu6 & Agyhu6);
assign Mmyhu6 = (Ru3iu6 & Xj3iu6);
assign Ru3iu6 = (~(Yu3iu6 & Fv3iu6));
assign Fv3iu6 = (Mv3iu6 & Tv3iu6);
assign Tv3iu6 = (Aw3iu6 | N73iu6);
assign N73iu6 = (~(Hw3iu6 & P5zhu6));
assign P5zhu6 = (!Ulnhu6);
assign Hw3iu6 = (~(Pyyhu6 & Mdhpw6[0]));
assign Pyyhu6 = (~(Qgzhu6 | O8zhu6));
assign Qgzhu6 = (!Mdhpw6[2]);
assign Mv3iu6 = (Ow3iu6 & P13iu6);
assign P13iu6 = (!Vmdpw6);
assign Yu3iu6 = (Rgnhu6 & Z63iu6);
assign Du3iu6 = (Xj3iu6 ? Vw3iu6 : A1zhu6);
assign Vw3iu6 = (T0zhu6 & Rzyhu6);
assign A1zhu6 = (~(Y7yhu6 | Ighpw6[0]));
assign It3iu6 = (Hknhu6 ? Jx3iu6 : Cx3iu6);
assign Jx3iu6 = (Ey3iu6 ? Xx3iu6 : Qx3iu6);
assign Qx3iu6 = (U5yhu6 & Ly3iu6);
assign Ly3iu6 = (~(Sy3iu6 & Zy3iu6));
assign Zy3iu6 = (Gz3iu6 & Y7yhu6);
assign Y7yhu6 = (~(Nz3iu6 & Ighpw6[2]));
assign Nz3iu6 = (~(Wdyhu6 | Ighpw6[1]));
assign Gz3iu6 = (~(T0zhu6 | Agyhu6));
assign T0zhu6 = (Gjyhu6 & Vuyhu6);
assign Sy3iu6 = (Uz3iu6 & B04iu6);
assign B04iu6 = (C9zhu6 | Vmzhu6);
assign Uz3iu6 = (I04iu6 & Joyhu6);
assign Joyhu6 = (~(P04iu6 & Epyhu6));
assign P04iu6 = (~(Deyhu6 | Ighpw6[2]));
assign I04iu6 = (~(Gjyhu6 & Eiyhu6));
assign Gjyhu6 = (~(C9zhu6 | Wdyhu6));
assign C9zhu6 = (!Cvyhu6);
assign Cx3iu6 = (~(Ey3iu6 & Xx3iu6));
assign Xx3iu6 = (~(W04iu6 & D14iu6));
assign D14iu6 = (~(K14iu6 & Z4yhu6));
assign K14iu6 = (Mdhpw6[0] & SWDO);
assign W04iu6 = (~(Mdhpw6[3] & R14iu6));
assign R14iu6 = (L02iu6 | R7yhu6);
assign R7yhu6 = (!Mdhpw6[0]);
assign L02iu6 = (!Z4yhu6);
assign Ey3iu6 = (Y14iu6 | Z4yhu6);
assign Z4yhu6 = (Ighpw6[5] & Vx2iu6);
assign Kfxhu6 = (M24iu6 ? F24iu6 : Aphpw6[1]);
assign F24iu6 = (T24iu6 & A34iu6);
assign Dfxhu6 = (M24iu6 ? H34iu6 : Cynhu6);
assign Wexhu6 = (M24iu6 ? O34iu6 : Aphpw6[2]);
assign M24iu6 = (V34iu6 & C44iu6);
assign Pexhu6 = (Sm1iu6 ? J44iu6 : Jshpw6[10]);
assign Iexhu6 = (Sm1iu6 ? Q44iu6 : Jshpw6[11]);
assign Bexhu6 = (Sm1iu6 ? X44iu6 : Jshpw6[12]);
assign Udxhu6 = (Sm1iu6 ? E54iu6 : Jshpw6[13]);
assign Ndxhu6 = (Sm1iu6 ? L54iu6 : Jshpw6[14]);
assign Gdxhu6 = (Sm1iu6 ? S54iu6 : Jshpw6[15]);
assign Zcxhu6 = (Sm1iu6 ? Z54iu6 : Jshpw6[16]);
assign Scxhu6 = (Sm1iu6 ? G64iu6 : Jshpw6[17]);
assign Lcxhu6 = (Sm1iu6 ? N64iu6 : Jshpw6[18]);
assign Ecxhu6 = (Sm1iu6 ? U64iu6 : Jshpw6[19]);
assign Xbxhu6 = (Sm1iu6 ? B74iu6 : Jshpw6[20]);
assign Qbxhu6 = (Sm1iu6 ? I74iu6 : Jshpw6[21]);
assign Jbxhu6 = (Sm1iu6 ? P74iu6 : Jshpw6[22]);
assign Cbxhu6 = (Sm1iu6 ? W74iu6 : Jshpw6[23]);
assign Vaxhu6 = (Sm1iu6 ? D84iu6 : Jshpw6[24]);
assign Oaxhu6 = (Sm1iu6 ? K84iu6 : Jshpw6[25]);
assign Haxhu6 = (Sm1iu6 ? R84iu6 : Jshpw6[26]);
assign Aaxhu6 = (Sm1iu6 ? Y84iu6 : Jshpw6[27]);
assign T9xhu6 = (Sm1iu6 ? F94iu6 : Jshpw6[28]);
assign M9xhu6 = (Sm1iu6 ? M94iu6 : Jshpw6[29]);
assign F9xhu6 = (Sm1iu6 ? T94iu6 : Jshpw6[30]);
assign Y8xhu6 = (~(Aa4iu6 & Ha4iu6));
assign Ha4iu6 = (~(Gmhpw6[0] & Oa4iu6));
assign Aa4iu6 = (Va4iu6 & Cb4iu6);
assign Cb4iu6 = (~(T24iu6 & Sm1iu6));
assign Va4iu6 = (~(Tnhpw6[0] & Jb4iu6));
assign R8xhu6 = (~(Qb4iu6 & Xb4iu6));
assign Xb4iu6 = (~(Gmhpw6[1] & Oa4iu6));
assign Qb4iu6 = (Ec4iu6 & Lc4iu6);
assign Lc4iu6 = (~(Sm1iu6 & O34iu6));
assign Ec4iu6 = (~(Tnhpw6[1] & Jb4iu6));
assign K8xhu6 = (~(Sc4iu6 & Zc4iu6));
assign Zc4iu6 = (~(Gmhpw6[2] & Oa4iu6));
assign Sc4iu6 = (Gd4iu6 & Nd4iu6);
assign Nd4iu6 = (~(Ud4iu6 & Sm1iu6));
assign Gd4iu6 = (~(Tnhpw6[2] & Jb4iu6));
assign D8xhu6 = (~(Be4iu6 & Ie4iu6));
assign Ie4iu6 = (~(Gmhpw6[3] & Oa4iu6));
assign Be4iu6 = (Pe4iu6 & We4iu6);
assign We4iu6 = (~(Df4iu6 & Sm1iu6));
assign Pe4iu6 = (~(Tnhpw6[3] & Jb4iu6));
assign W7xhu6 = (~(Kf4iu6 & Rf4iu6));
assign Rf4iu6 = (~(Gmhpw6[4] & Oa4iu6));
assign Kf4iu6 = (Yf4iu6 & Fg4iu6);
assign Fg4iu6 = (~(H34iu6 & Sm1iu6));
assign Yf4iu6 = (~(Jshpw6[4] & Jb4iu6));
assign P7xhu6 = (~(Mg4iu6 & Tg4iu6));
assign Tg4iu6 = (~(Gmhpw6[5] & Oa4iu6));
assign Mg4iu6 = (Ah4iu6 & Hh4iu6);
assign Hh4iu6 = (~(Oh4iu6 & Sm1iu6));
assign Ah4iu6 = (~(Jshpw6[5] & Jb4iu6));
assign I7xhu6 = (~(Vh4iu6 & Ci4iu6));
assign Ci4iu6 = (~(Gmhpw6[6] & Oa4iu6));
assign Vh4iu6 = (Ji4iu6 & Qi4iu6);
assign Qi4iu6 = (~(Xi4iu6 & Sm1iu6));
assign Ji4iu6 = (~(Jshpw6[6] & Jb4iu6));
assign B7xhu6 = (~(Ej4iu6 & Lj4iu6));
assign Lj4iu6 = (~(Gmhpw6[7] & Oa4iu6));
assign Ej4iu6 = (Sj4iu6 & Zj4iu6);
assign Zj4iu6 = (~(Gk4iu6 & Sm1iu6));
assign Sj4iu6 = (~(Jshpw6[7] & Jb4iu6));
assign U6xhu6 = (~(Nk4iu6 & Uk4iu6));
assign Uk4iu6 = (~(Gmhpw6[8] & Oa4iu6));
assign Nk4iu6 = (Bl4iu6 & Il4iu6);
assign Il4iu6 = (~(Sm1iu6 & Pl4iu6));
assign Bl4iu6 = (~(Jshpw6[8] & Jb4iu6));
assign N6xhu6 = (~(Wl4iu6 & Dm4iu6));
assign Dm4iu6 = (~(Gmhpw6[9] & Oa4iu6));
assign Wl4iu6 = (Km4iu6 & Rm4iu6);
assign Rm4iu6 = (~(Sm1iu6 & Ym4iu6));
assign Sm1iu6 = (~(Jb4iu6 | Oa4iu6));
assign Km4iu6 = (~(Jshpw6[9] & Jb4iu6));
assign Jb4iu6 = (~(Fn4iu6 | Oa4iu6));
assign Oa4iu6 = (Mn4iu6 & Tn4iu6);
assign Tn4iu6 = (Ao4iu6 & Pqzhu6);
assign Ao4iu6 = (~(Lf1iu6 | Ho4iu6));
assign Lf1iu6 = (HRESP & R0nhu6);
assign Mn4iu6 = (Cynhu6 & Tszhu6);
assign Tszhu6 = (Oo4iu6 & Sqhpw6[1]);
assign Oo4iu6 = (~(Fszhu6 | Sqhpw6[0]));
assign Fn4iu6 = (V34iu6 & Vo4iu6);
assign V34iu6 = (Cp4iu6 & Jp4iu6);
assign Jp4iu6 = (Qp4iu6 & Xp4iu6);
assign Qp4iu6 = (~(Ho4iu6 | Eq4iu6));
assign Cp4iu6 = (Lq4iu6 & Sqhpw6[1]);
assign Lq4iu6 = (~(Gpzhu6 | Sq4iu6));
assign G6xhu6 = (!Zq4iu6);
assign Zq4iu6 = (Nr4iu6 ? Sq4iu6 : Gr4iu6);
assign Gr4iu6 = (~(A2nhu6 & Ur4iu6));
assign Z5xhu6 = (Bs4iu6 ? Lwgpw6[0] : T24iu6);
assign S5xhu6 = (Bs4iu6 ? Lwgpw6[2] : Ud4iu6);
assign L5xhu6 = (Bs4iu6 ? Lwgpw6[1] : O34iu6);
assign Bs4iu6 = (Is4iu6 | Ps4iu6);
assign Is4iu6 = (!Ws4iu6);
assign E5xhu6 = (Kt4iu6 ? Dt4iu6 : Vchhu6);
assign Kt4iu6 = (HREADY & Rt4iu6);
assign Rt4iu6 = (~(Yt4iu6 & Fu4iu6));
assign Fu4iu6 = (~(Mu4iu6 | Tu4iu6));
assign Yt4iu6 = (~(Dt4iu6 | Av4iu6));
assign Av4iu6 = (~(Hv4iu6 | DBGRESTART));
assign Dt4iu6 = (~(Ov4iu6 & Vv4iu6));
assign Vv4iu6 = (Cw4iu6 & Jw4iu6);
assign Cw4iu6 = (Qw4iu6 & Xw4iu6);
assign Ov4iu6 = (~(Ex4iu6 | Lx4iu6));
assign X4xhu6 = (~(Sx4iu6 & Zx4iu6));
assign Zx4iu6 = (Gy4iu6 & Ny4iu6);
assign Ny4iu6 = (~(Hrfpw6[16] & Uy4iu6));
assign Gy4iu6 = (Bz4iu6 & Iz4iu6);
assign Bz4iu6 = (~(Pz4iu6 & Wz4iu6));
assign Sx4iu6 = (D05iu6 & K05iu6);
assign K05iu6 = (~(R05iu6 & S1ehu6));
assign D05iu6 = (Y05iu6 & F15iu6);
assign F15iu6 = (~(M15iu6 & T15iu6));
assign Y05iu6 = (~(Ppfpw6[16] & A25iu6));
assign Q4xhu6 = (O25iu6 ? X3fpw6[1] : H25iu6);
assign H25iu6 = (~(V25iu6 & C35iu6));
assign C35iu6 = (J35iu6 & Q35iu6);
assign Q35iu6 = (X35iu6 & E45iu6);
assign X35iu6 = (~(L45iu6 & S45iu6));
assign S45iu6 = (~(Z45iu6 & G55iu6));
assign Z45iu6 = (B65iu6 ? U55iu6 : N55iu6);
assign U55iu6 = (~(I65iu6 & P65iu6));
assign J35iu6 = (W65iu6 & D75iu6);
assign D75iu6 = (~(D7fpw6[4] & K75iu6));
assign W65iu6 = (R75iu6 | P65iu6);
assign V25iu6 = (Y75iu6 & F85iu6);
assign Y75iu6 = (M85iu6 & T85iu6);
assign T85iu6 = (~(A95iu6 & D7fpw6[1]));
assign M85iu6 = (H95iu6 | O95iu6);
assign J4xhu6 = (Fsdhu6 ? Ca5iu6 : V95iu6);
assign Ca5iu6 = (~(Ja5iu6 & Qa5iu6));
assign V95iu6 = (~(Xa5iu6 & Eb5iu6));
assign Eb5iu6 = (Lb5iu6 & Sb5iu6);
assign Lb5iu6 = (~(RXEV | TXEV));
assign Xa5iu6 = (Zb5iu6 & Gc5iu6);
assign Zb5iu6 = (Nc5iu6 & Uc5iu6);
assign Nc5iu6 = (~(Gfghu6 & Bd5iu6));
assign Bd5iu6 = (~(Id5iu6 & Pd5iu6));
assign Pd5iu6 = (Wd5iu6 & De5iu6);
assign De5iu6 = (Ke5iu6 & Re5iu6);
assign Re5iu6 = (Ye5iu6 & Ff5iu6);
assign Ff5iu6 = (Mf5iu6 & Tf5iu6);
assign Tf5iu6 = (Ag5iu6 | Yyghu6);
assign Mf5iu6 = (Hg5iu6 & Og5iu6);
assign Og5iu6 = (~(Vg5iu6 & Ch5iu6));
assign Vg5iu6 = (HWDATA[28] & Jh5iu6);
assign Hg5iu6 = (Qh5iu6 | Zlghu6);
assign Ye5iu6 = (Xh5iu6 & Ei5iu6);
assign Ei5iu6 = (Li5iu6 | Righu6);
assign Xh5iu6 = (~(Cyohu6 & Si5iu6));
assign Si5iu6 = (!Odgpw6[31]);
assign Ke5iu6 = (Zi5iu6 & Gj5iu6);
assign Gj5iu6 = (Nj5iu6 & Uj5iu6);
assign Uj5iu6 = (~(Xyohu6 & Bk5iu6));
assign Bk5iu6 = (!Odgpw6[28]);
assign Nj5iu6 = (Ik5iu6 & Pk5iu6);
assign Pk5iu6 = (~(Jyohu6 & Wk5iu6));
assign Wk5iu6 = (!Odgpw6[30]);
assign Ik5iu6 = (~(Qyohu6 & Dl5iu6));
assign Dl5iu6 = (!Odgpw6[29]);
assign Zi5iu6 = (Kl5iu6 & Rl5iu6);
assign Rl5iu6 = (~(Ezohu6 & Yl5iu6));
assign Yl5iu6 = (!Odgpw6[27]);
assign Kl5iu6 = (~(Lzohu6 & Fm5iu6));
assign Fm5iu6 = (!Odgpw6[26]);
assign Wd5iu6 = (Mm5iu6 & Tm5iu6);
assign Tm5iu6 = (An5iu6 & Hn5iu6);
assign Hn5iu6 = (On5iu6 & Vn5iu6);
assign Vn5iu6 = (~(G0phu6 & Co5iu6));
assign Co5iu6 = (!Odgpw6[21]);
assign On5iu6 = (Jo5iu6 & Qo5iu6);
assign Qo5iu6 = (~(Szohu6 & Xo5iu6));
assign Xo5iu6 = (!Odgpw6[23]);
assign Jo5iu6 = (~(Zzohu6 & Ep5iu6));
assign Ep5iu6 = (!Odgpw6[22]);
assign An5iu6 = (Lp5iu6 & Sp5iu6);
assign Sp5iu6 = (~(N0phu6 & Zp5iu6));
assign Zp5iu6 = (!Odgpw6[20]);
assign Lp5iu6 = (~(U0phu6 & Gq5iu6));
assign Gq5iu6 = (!Odgpw6[19]);
assign Mm5iu6 = (Nq5iu6 & Uq5iu6);
assign Uq5iu6 = (Br5iu6 & Ir5iu6);
assign Ir5iu6 = (~(B1phu6 & Pr5iu6));
assign Pr5iu6 = (!Odgpw6[18]);
assign Br5iu6 = (~(I1phu6 & Wr5iu6));
assign Wr5iu6 = (!Odgpw6[17]);
assign Nq5iu6 = (Ds5iu6 & Ks5iu6);
assign Ks5iu6 = (~(P1phu6 & Rs5iu6));
assign Rs5iu6 = (!Odgpw6[16]);
assign Ds5iu6 = (~(W1phu6 & Ys5iu6));
assign Ys5iu6 = (!Odgpw6[15]);
assign Id5iu6 = (Ft5iu6 & Mt5iu6);
assign Mt5iu6 = (Tt5iu6 & Au5iu6);
assign Au5iu6 = (Hu5iu6 & Ou5iu6);
assign Ou5iu6 = (Vu5iu6 & Cv5iu6);
assign Cv5iu6 = (~(R2phu6 & Jv5iu6));
assign Jv5iu6 = (!Odgpw6[12]);
assign Vu5iu6 = (Qv5iu6 & Xv5iu6);
assign Xv5iu6 = (~(D2phu6 & Ew5iu6));
assign Ew5iu6 = (!Odgpw6[14]);
assign Qv5iu6 = (~(K2phu6 & Lw5iu6));
assign Lw5iu6 = (!Odgpw6[13]);
assign Hu5iu6 = (Sw5iu6 & Zw5iu6);
assign Zw5iu6 = (~(Y2phu6 & Gx5iu6));
assign Gx5iu6 = (!Odgpw6[11]);
assign Sw5iu6 = (~(F3phu6 & Nx5iu6));
assign Nx5iu6 = (!Odgpw6[10]);
assign Tt5iu6 = (Ux5iu6 & By5iu6);
assign By5iu6 = (Iy5iu6 & Py5iu6);
assign Py5iu6 = (~(M3phu6 & Wy5iu6));
assign Wy5iu6 = (!Odgpw6[7]);
assign Iy5iu6 = (~(T3phu6 & Dz5iu6));
assign Dz5iu6 = (!Odgpw6[6]);
assign Ux5iu6 = (Kz5iu6 & Rz5iu6);
assign Rz5iu6 = (~(A4phu6 & Yz5iu6));
assign Yz5iu6 = (!Odgpw6[5]);
assign Kz5iu6 = (~(H4phu6 & F06iu6));
assign F06iu6 = (!Odgpw6[4]);
assign Ft5iu6 = (M06iu6 & T06iu6);
assign T06iu6 = (A16iu6 & H16iu6);
assign H16iu6 = (O16iu6 & V16iu6);
assign V16iu6 = (~(C5phu6 & C26iu6));
assign C26iu6 = (!Odgpw6[1]);
assign O16iu6 = (J26iu6 & Q26iu6);
assign Q26iu6 = (~(O4phu6 & X26iu6));
assign X26iu6 = (!Odgpw6[3]);
assign J26iu6 = (~(V4phu6 & E36iu6));
assign E36iu6 = (!Odgpw6[2]);
assign A16iu6 = (L36iu6 & S36iu6);
assign S36iu6 = (~(J5phu6 & Z36iu6));
assign Z36iu6 = (!Odgpw6[0]);
assign L36iu6 = (~(Bxdpw6 & G46iu6));
assign G46iu6 = (!Odgpw6[8]);
assign Bxdpw6 = (N46iu6 & U46iu6);
assign U46iu6 = (~(B56iu6 & I56iu6));
assign I56iu6 = (~(Sodpw6 & IRQ[8]));
assign B56iu6 = (P56iu6 & W56iu6);
assign P56iu6 = (~(Odgpw6[8] & D66iu6));
assign D66iu6 = (~(K66iu6 & HWDATA[8]));
assign M06iu6 = (R66iu6 & Y66iu6);
assign Y66iu6 = (F76iu6 & M76iu6);
assign M76iu6 = (~(Uwdpw6 & T76iu6));
assign T76iu6 = (!Odgpw6[9]);
assign Uwdpw6 = (A86iu6 & H86iu6);
assign H86iu6 = (~(O86iu6 & V86iu6));
assign V86iu6 = (~(Cndpw6 & IRQ[9]));
assign O86iu6 = (C96iu6 & J96iu6);
assign C96iu6 = (~(Odgpw6[9] & Q96iu6));
assign Q96iu6 = (~(K66iu6 & HWDATA[9]));
assign F76iu6 = (~(Nwdpw6 & X96iu6));
assign X96iu6 = (!Odgpw6[24]);
assign Nwdpw6 = (Ea6iu6 & La6iu6);
assign La6iu6 = (~(Sa6iu6 & Za6iu6));
assign Za6iu6 = (~(Wqdpw6 & IRQ[24]));
assign Sa6iu6 = (Gb6iu6 & Nb6iu6);
assign Gb6iu6 = (~(Odgpw6[24] & Ub6iu6));
assign Ub6iu6 = (~(K66iu6 & HWDATA[24]));
assign R66iu6 = (Bc6iu6 & Ic6iu6);
assign Ic6iu6 = (~(Gwdpw6 & Pc6iu6));
assign Pc6iu6 = (!Odgpw6[25]);
assign Gwdpw6 = (Wc6iu6 & Dd6iu6);
assign Dd6iu6 = (~(Kd6iu6 & Rd6iu6));
assign Rd6iu6 = (~(Krdpw6 & IRQ[25]));
assign Kd6iu6 = (Yd6iu6 & Fe6iu6);
assign Yd6iu6 = (~(Odgpw6[25] & Me6iu6));
assign Me6iu6 = (~(K66iu6 & HWDATA[25]));
assign Bc6iu6 = (~(Npghu6 & Te6iu6));
assign Npghu6 = (Af6iu6 & Hf6iu6);
assign Hf6iu6 = (~(Of6iu6 & Vf6iu6));
assign Vf6iu6 = (~(Evdpw6 & NMI));
assign Of6iu6 = (Cg6iu6 & Jg6iu6);
assign Cg6iu6 = (Te6iu6 | Qg6iu6);
assign C4xhu6 = (Eh6iu6 ? R0nhu6 : Xg6iu6);
assign O3xhu6 = (~(Lh6iu6 & Sh6iu6));
assign Sh6iu6 = (Zh6iu6 | HREADY);
assign Lh6iu6 = (Gi6iu6 & Ni6iu6);
assign Gi6iu6 = (~(Ui6iu6 & Nr4iu6));
assign Ui6iu6 = (~(Bj6iu6 ^ Jshpw6[5]));
assign H3xhu6 = (~(Ij6iu6 & Pj6iu6));
assign Pj6iu6 = (Wj6iu6 | HREADY);
assign Ij6iu6 = (Dk6iu6 & Ni6iu6);
assign Dk6iu6 = (~(Kk6iu6 & Nr4iu6));
assign Kk6iu6 = (~(Bj6iu6 ^ Jshpw6[13]));
assign A3xhu6 = (~(Rk6iu6 & Yk6iu6));
assign Yk6iu6 = (Fl6iu6 | HREADY);
assign Rk6iu6 = (Ml6iu6 & Ni6iu6);
assign Ml6iu6 = (~(Tl6iu6 & Nr4iu6));
assign Tl6iu6 = (~(Am6iu6 ^ Jshpw6[4]));
assign T2xhu6 = (~(Hm6iu6 & Om6iu6));
assign Om6iu6 = (Vm6iu6 | HREADY);
assign Hm6iu6 = (Cn6iu6 & Ni6iu6);
assign Cn6iu6 = (~(Jn6iu6 & Nr4iu6));
assign Jn6iu6 = (~(Am6iu6 ^ Jshpw6[12]));
assign M2xhu6 = (~(Qn6iu6 & Xn6iu6));
assign Xn6iu6 = (Eo6iu6 | HREADY);
assign Qn6iu6 = (Lo6iu6 & Ni6iu6);
assign Lo6iu6 = (~(Nr4iu6 & So6iu6));
assign So6iu6 = (~(Zo6iu6 ^ Jshpw6[15]));
assign F2xhu6 = (~(Gp6iu6 & Np6iu6));
assign Np6iu6 = (~(X8hpw6[1] & Eh6iu6));
assign Gp6iu6 = (Up6iu6 & Ni6iu6);
assign Up6iu6 = (Bq6iu6 | Iq6iu6);
assign Y1xhu6 = (~(Pq6iu6 & Wq6iu6));
assign Wq6iu6 = (Dr6iu6 | HREADY);
assign Pq6iu6 = (Kr6iu6 & Ni6iu6);
assign Ni6iu6 = (~(Nr4iu6 & Rr6iu6));
assign Rr6iu6 = (~(Yr6iu6 & Fs6iu6));
assign Yr6iu6 = (Ms6iu6 & Ts6iu6);
assign Ts6iu6 = (At6iu6 & Ht6iu6);
assign Ht6iu6 = (Wqzhu6 | Aphpw6[2]);
assign Ms6iu6 = (Ot6iu6 & Vt6iu6);
assign Vt6iu6 = (Cu6iu6 | Jshpw6[8]);
assign Cu6iu6 = (!Jshpw6[11]);
assign Ot6iu6 = (Jshpw6[10] ? Qu6iu6 : Ju6iu6);
assign Qu6iu6 = (Jshpw6[11] & Xu6iu6);
assign Xu6iu6 = (~(Ev6iu6 & Lv6iu6));
assign Lv6iu6 = (~(Sv6iu6 & Zv6iu6));
assign Zv6iu6 = (Gw6iu6 & Nw6iu6);
assign Gw6iu6 = (Uw6iu6 & Bx6iu6);
assign Sv6iu6 = (Ix6iu6 & Px6iu6);
assign Px6iu6 = (Jshpw6[6] ? Dy6iu6 : Wx6iu6);
assign Dy6iu6 = (~(Ky6iu6 | Ry6iu6));
assign Wx6iu6 = (Yy6iu6 & Bj6iu6);
assign Yy6iu6 = (~(Jshpw6[7] | Jshpw6[9]));
assign Ix6iu6 = (Fz6iu6 & Mz6iu6);
assign Fz6iu6 = (~(Jshpw6[4] ^ Jshpw6[5]));
assign Ev6iu6 = (~(Tz6iu6 & A07iu6));
assign A07iu6 = (Jshpw6[6] & H07iu6);
assign H07iu6 = (~(O07iu6 & V07iu6));
assign V07iu6 = (~(C17iu6 & J17iu6));
assign C17iu6 = (~(Am6iu6 | Bj6iu6));
assign O07iu6 = (~(Q17iu6 & X17iu6));
assign X17iu6 = (~(E27iu6 & L27iu6));
assign E27iu6 = (~(S27iu6 & Z27iu6));
assign S27iu6 = (Bx6iu6 ? Jshpw6[13] : G37iu6);
assign Q17iu6 = (~(N37iu6 & U37iu6));
assign N37iu6 = (~(B47iu6 & Jshpw6[4]));
assign B47iu6 = (~(I47iu6 | P47iu6));
assign Tz6iu6 = (~(Iq6iu6 | Ky6iu6));
assign Iq6iu6 = (!Jshpw6[9]);
assign Ju6iu6 = (W47iu6 & D57iu6);
assign D57iu6 = (K57iu6 & Ky6iu6);
assign Ky6iu6 = (!Jshpw6[7]);
assign K57iu6 = (~(Jshpw6[8] | Jshpw6[9]));
assign W47iu6 = (R57iu6 & Zo6iu6);
assign Zo6iu6 = (!Jshpw6[6]);
assign R57iu6 = (~(Y57iu6 & F67iu6));
assign F67iu6 = (~(M67iu6 & T67iu6));
assign T67iu6 = (A77iu6 & Mz6iu6);
assign A77iu6 = (~(Bx6iu6 | Jshpw6[15]));
assign M67iu6 = (H77iu6 & G37iu6);
assign G37iu6 = (~(Jshpw6[14] | Jshpw6[13]));
assign H77iu6 = (Jshpw6[5] ? V77iu6 : O77iu6);
assign V77iu6 = (Am6iu6 | Bj6iu6);
assign O77iu6 = (C87iu6 & J87iu6);
assign J87iu6 = (Bj6iu6 | Jshpw6[4]);
assign C87iu6 = (I47iu6 ? P47iu6 : Ry6iu6);
assign Ry6iu6 = (!Jshpw6[4]);
assign Y57iu6 = (~(U37iu6 & Q87iu6));
assign Q87iu6 = (J17iu6 | X87iu6);
assign X87iu6 = (E97iu6 & L97iu6);
assign L97iu6 = (S97iu6 & Jshpw6[13]);
assign S97iu6 = (Z97iu6 & Bx6iu6);
assign Z97iu6 = (~(Jshpw6[14] & Uw6iu6));
assign Uw6iu6 = (Am6iu6 | P47iu6);
assign Am6iu6 = (!I47iu6);
assign E97iu6 = (~(Ga7iu6 | Na7iu6));
assign Na7iu6 = (!Z27iu6);
assign Z27iu6 = (Ua7iu6 & Mz6iu6);
assign Ua7iu6 = (~(Jshpw6[14] ^ Jshpw6[15]));
assign Ga7iu6 = (Jshpw6[4] ? I47iu6 : Bb7iu6);
assign Bb7iu6 = (~(I47iu6 | Bj6iu6));
assign Bj6iu6 = (!P47iu6);
assign J17iu6 = (~(L27iu6 | Jshpw6[4]));
assign L27iu6 = (~(Ib7iu6 & Pb7iu6));
assign Pb7iu6 = (Wb7iu6 & Jshpw6[17]);
assign Wb7iu6 = (Jshpw6[16] & Jshpw6[12]);
assign Ib7iu6 = (Dc7iu6 & Nw6iu6);
assign Nw6iu6 = (Kc7iu6 & Jshpw6[15]);
assign Dc7iu6 = (Jshpw6[19] & Jshpw6[18]);
assign U37iu6 = (!Jshpw6[5]);
assign Nr4iu6 = (!Bq6iu6);
assign Kr6iu6 = (Bq6iu6 | Bx6iu6);
assign R1xhu6 = (Rc7iu6 ? E5hhu6 : D84iu6);
assign K1xhu6 = (Rc7iu6 ? H2hhu6 : T24iu6);
assign D1xhu6 = (Rc7iu6 ? S3hhu6 : J44iu6);
assign Rc7iu6 = (~(Yc7iu6 & A2nhu6));
assign W0xhu6 = (Fd7iu6 ? Jehhu6 : T24iu6);
assign P0xhu6 = (Fd7iu6 ? Hbhhu6 : Ud4iu6);
assign Fd7iu6 = (!Tu4iu6);
assign I0xhu6 = (Tu4iu6 ? Df4iu6 : P9hhu6);
assign B0xhu6 = (Md7iu6 ? Togpw6[2] : Ud4iu6);
assign Uzwhu6 = (Md7iu6 ? Ligpw6[28] : Lm1iu6);
assign Nzwhu6 = (Md7iu6 ? Ligpw6[27] : T94iu6);
assign Gzwhu6 = (Md7iu6 ? Togpw6[28] : F94iu6);
assign Zywhu6 = (Md7iu6 ? Togpw6[27] : Y84iu6);
assign Sywhu6 = (Md7iu6 ? Togpw6[26] : R84iu6);
assign Lywhu6 = (Md7iu6 ? Togpw6[25] : K84iu6);
assign Eywhu6 = (Md7iu6 ? Togpw6[24] : D84iu6);
assign Xxwhu6 = (Md7iu6 ? Togpw6[23] : W74iu6);
assign Qxwhu6 = (Md7iu6 ? Togpw6[22] : P74iu6);
assign Jxwhu6 = (Md7iu6 ? Togpw6[21] : I74iu6);
assign Cxwhu6 = (Md7iu6 ? Togpw6[20] : B74iu6);
assign Vwwhu6 = (Md7iu6 ? Togpw6[19] : U64iu6);
assign Owwhu6 = (Md7iu6 ? Togpw6[18] : N64iu6);
assign Hwwhu6 = (Md7iu6 ? Togpw6[17] : G64iu6);
assign Awwhu6 = (Md7iu6 ? Togpw6[16] : Z54iu6);
assign Tvwhu6 = (Md7iu6 ? Togpw6[15] : S54iu6);
assign Mvwhu6 = (Md7iu6 ? Togpw6[14] : L54iu6);
assign Fvwhu6 = (Md7iu6 ? Togpw6[13] : E54iu6);
assign Yuwhu6 = (Md7iu6 ? Togpw6[12] : X44iu6);
assign Ruwhu6 = (Md7iu6 ? Togpw6[11] : Q44iu6);
assign Kuwhu6 = (Md7iu6 ? Togpw6[10] : J44iu6);
assign Duwhu6 = (Md7iu6 ? Togpw6[9] : Ym4iu6);
assign Wtwhu6 = (Md7iu6 ? Togpw6[8] : Pl4iu6);
assign Ptwhu6 = (Md7iu6 ? Togpw6[7] : Gk4iu6);
assign Itwhu6 = (Md7iu6 ? Togpw6[6] : Xi4iu6);
assign Btwhu6 = (Md7iu6 ? Togpw6[5] : Oh4iu6);
assign Uswhu6 = (Md7iu6 ? Togpw6[4] : H34iu6);
assign Nswhu6 = (Md7iu6 ? Togpw6[3] : Df4iu6);
assign Gswhu6 = (Md7iu6 ? Qhhhu6 : T24iu6);
assign Md7iu6 = (~(A2nhu6 & Vr1iu6));
assign Zrwhu6 = (Td7iu6 ? Gqgpw6[2] : Ud4iu6);
assign Srwhu6 = (Td7iu6 ? Akgpw6[28] : Lm1iu6);
assign Lrwhu6 = (Td7iu6 ? Akgpw6[27] : T94iu6);
assign Erwhu6 = (Td7iu6 ? Gqgpw6[28] : F94iu6);
assign Xqwhu6 = (Td7iu6 ? Gqgpw6[27] : Y84iu6);
assign Qqwhu6 = (Td7iu6 ? Gqgpw6[26] : R84iu6);
assign Jqwhu6 = (Td7iu6 ? Gqgpw6[25] : K84iu6);
assign Cqwhu6 = (Td7iu6 ? Gqgpw6[24] : D84iu6);
assign Vpwhu6 = (Td7iu6 ? Gqgpw6[23] : W74iu6);
assign Opwhu6 = (Td7iu6 ? Gqgpw6[22] : P74iu6);
assign Hpwhu6 = (Td7iu6 ? Gqgpw6[21] : I74iu6);
assign Apwhu6 = (Td7iu6 ? Gqgpw6[20] : B74iu6);
assign Towhu6 = (Td7iu6 ? Gqgpw6[19] : U64iu6);
assign Mowhu6 = (Td7iu6 ? Gqgpw6[18] : N64iu6);
assign Fowhu6 = (Td7iu6 ? Gqgpw6[17] : G64iu6);
assign Ynwhu6 = (Td7iu6 ? Gqgpw6[16] : Z54iu6);
assign Rnwhu6 = (Td7iu6 ? Gqgpw6[15] : S54iu6);
assign Knwhu6 = (Td7iu6 ? Gqgpw6[14] : L54iu6);
assign Dnwhu6 = (Td7iu6 ? Gqgpw6[13] : E54iu6);
assign Wmwhu6 = (Td7iu6 ? Gqgpw6[12] : X44iu6);
assign Pmwhu6 = (Td7iu6 ? Gqgpw6[11] : Q44iu6);
assign Imwhu6 = (Td7iu6 ? Gqgpw6[10] : J44iu6);
assign Bmwhu6 = (Td7iu6 ? Gqgpw6[9] : Ym4iu6);
assign Ulwhu6 = (Td7iu6 ? Gqgpw6[8] : Pl4iu6);
assign Nlwhu6 = (Td7iu6 ? Gqgpw6[7] : Gk4iu6);
assign Glwhu6 = (Td7iu6 ? Gqgpw6[6] : Xi4iu6);
assign Zkwhu6 = (Td7iu6 ? Gqgpw6[5] : Oh4iu6);
assign Skwhu6 = (Td7iu6 ? Gqgpw6[4] : H34iu6);
assign Lkwhu6 = (Td7iu6 ? Gqgpw6[3] : Df4iu6);
assign Ekwhu6 = (Td7iu6 ? Ijhhu6 : T24iu6);
assign Td7iu6 = (~(A2nhu6 & Xs1iu6));
assign Xjwhu6 = (Ae7iu6 ? Trgpw6[2] : Ud4iu6);
assign Qjwhu6 = (Ae7iu6 ? Plgpw6[28] : Lm1iu6);
assign Jjwhu6 = (Ae7iu6 ? Plgpw6[27] : T94iu6);
assign Cjwhu6 = (Ae7iu6 ? Trgpw6[28] : F94iu6);
assign Viwhu6 = (Ae7iu6 ? Trgpw6[27] : Y84iu6);
assign Oiwhu6 = (Ae7iu6 ? Trgpw6[26] : R84iu6);
assign Hiwhu6 = (Ae7iu6 ? Trgpw6[25] : K84iu6);
assign Aiwhu6 = (Ae7iu6 ? Trgpw6[24] : D84iu6);
assign Thwhu6 = (Ae7iu6 ? Trgpw6[23] : W74iu6);
assign Mhwhu6 = (Ae7iu6 ? Trgpw6[22] : P74iu6);
assign Fhwhu6 = (Ae7iu6 ? Trgpw6[21] : I74iu6);
assign Ygwhu6 = (Ae7iu6 ? Trgpw6[20] : B74iu6);
assign Rgwhu6 = (Ae7iu6 ? Trgpw6[19] : U64iu6);
assign Kgwhu6 = (Ae7iu6 ? Trgpw6[18] : N64iu6);
assign Dgwhu6 = (Ae7iu6 ? Trgpw6[17] : G64iu6);
assign Wfwhu6 = (Ae7iu6 ? Trgpw6[16] : Z54iu6);
assign Pfwhu6 = (Ae7iu6 ? Trgpw6[15] : S54iu6);
assign Ifwhu6 = (Ae7iu6 ? Trgpw6[14] : L54iu6);
assign Bfwhu6 = (Ae7iu6 ? Trgpw6[13] : E54iu6);
assign Uewhu6 = (Ae7iu6 ? Trgpw6[12] : X44iu6);
assign Newhu6 = (Ae7iu6 ? Trgpw6[11] : Q44iu6);
assign Gewhu6 = (Ae7iu6 ? Trgpw6[10] : J44iu6);
assign Zdwhu6 = (Ae7iu6 ? Trgpw6[9] : Ym4iu6);
assign Sdwhu6 = (Ae7iu6 ? Trgpw6[8] : Pl4iu6);
assign Ldwhu6 = (Ae7iu6 ? Trgpw6[7] : Gk4iu6);
assign Edwhu6 = (Ae7iu6 ? Trgpw6[6] : Xi4iu6);
assign Xcwhu6 = (Ae7iu6 ? Trgpw6[5] : Oh4iu6);
assign Qcwhu6 = (Ae7iu6 ? Trgpw6[4] : H34iu6);
assign Jcwhu6 = (Ae7iu6 ? Trgpw6[3] : Df4iu6);
assign Ccwhu6 = (Ae7iu6 ? Alhhu6 : T24iu6);
assign Ae7iu6 = (~(A2nhu6 & Dw1iu6));
assign Vbwhu6 = (He7iu6 ? Gtgpw6[2] : Ud4iu6);
assign Obwhu6 = (He7iu6 ? Engpw6[28] : Lm1iu6);
assign Hbwhu6 = (He7iu6 ? Engpw6[27] : T94iu6);
assign Abwhu6 = (He7iu6 ? Gtgpw6[28] : F94iu6);
assign Tawhu6 = (He7iu6 ? Gtgpw6[27] : Y84iu6);
assign Mawhu6 = (He7iu6 ? Gtgpw6[26] : R84iu6);
assign Fawhu6 = (He7iu6 ? Gtgpw6[25] : K84iu6);
assign Y9whu6 = (He7iu6 ? Gtgpw6[24] : D84iu6);
assign R9whu6 = (He7iu6 ? Gtgpw6[23] : W74iu6);
assign K9whu6 = (He7iu6 ? Gtgpw6[22] : P74iu6);
assign D9whu6 = (He7iu6 ? Gtgpw6[21] : I74iu6);
assign W8whu6 = (He7iu6 ? Gtgpw6[20] : B74iu6);
assign P8whu6 = (He7iu6 ? Gtgpw6[19] : U64iu6);
assign I8whu6 = (He7iu6 ? Gtgpw6[18] : N64iu6);
assign B8whu6 = (He7iu6 ? Gtgpw6[17] : G64iu6);
assign U7whu6 = (He7iu6 ? Gtgpw6[16] : Z54iu6);
assign N7whu6 = (He7iu6 ? Gtgpw6[15] : S54iu6);
assign G7whu6 = (He7iu6 ? Gtgpw6[14] : L54iu6);
assign Z6whu6 = (He7iu6 ? Gtgpw6[13] : E54iu6);
assign S6whu6 = (He7iu6 ? Gtgpw6[12] : X44iu6);
assign L6whu6 = (He7iu6 ? Gtgpw6[11] : Q44iu6);
assign E6whu6 = (He7iu6 ? Gtgpw6[10] : J44iu6);
assign X5whu6 = (He7iu6 ? Gtgpw6[9] : Ym4iu6);
assign Q5whu6 = (He7iu6 ? Gtgpw6[8] : Pl4iu6);
assign J5whu6 = (He7iu6 ? Gtgpw6[7] : Gk4iu6);
assign C5whu6 = (He7iu6 ? Gtgpw6[6] : Xi4iu6);
assign V4whu6 = (He7iu6 ? Gtgpw6[5] : Oh4iu6);
assign O4whu6 = (He7iu6 ? Gtgpw6[4] : H34iu6);
assign H4whu6 = (He7iu6 ? Gtgpw6[3] : Df4iu6);
assign A4whu6 = (He7iu6 ? Smhhu6 : T24iu6);
assign He7iu6 = (~(A2nhu6 & Cs1iu6));
assign T3whu6 = (Oe7iu6 ? T24iu6 : Kohhu6);
assign Oe7iu6 = (Ve7iu6 & A2nhu6);
assign M3whu6 = (Cf7iu6 ? Aygpw6[0] : T24iu6);
assign F3whu6 = (Cf7iu6 ? Aygpw6[4] : H34iu6);
assign Y2whu6 = (Cf7iu6 ? Aygpw6[3] : Df4iu6);
assign R2whu6 = (Cf7iu6 ? Aygpw6[2] : Ud4iu6);
assign K2whu6 = (Cf7iu6 ? Aygpw6[1] : O34iu6);
assign Cf7iu6 = (~(Jf7iu6 & A2nhu6));
assign D2whu6 = (Qf7iu6 ? Pzgpw6[0] : T24iu6);
assign W1whu6 = (Qf7iu6 ? E1hpw6[31] : Lm1iu6);
assign P1whu6 = (Qf7iu6 ? E1hpw6[30] : T94iu6);
assign I1whu6 = (Qf7iu6 ? E1hpw6[29] : M94iu6);
assign B1whu6 = (Qf7iu6 ? E1hpw6[28] : F94iu6);
assign U0whu6 = (Qf7iu6 ? E1hpw6[27] : Y84iu6);
assign N0whu6 = (Qf7iu6 ? E1hpw6[26] : R84iu6);
assign G0whu6 = (Qf7iu6 ? E1hpw6[25] : K84iu6);
assign Zzvhu6 = (Qf7iu6 ? E1hpw6[24] : D84iu6);
assign Szvhu6 = (Qf7iu6 ? E1hpw6[23] : W74iu6);
assign Lzvhu6 = (Qf7iu6 ? E1hpw6[22] : P74iu6);
assign Ezvhu6 = (Qf7iu6 ? E1hpw6[21] : I74iu6);
assign Xyvhu6 = (Qf7iu6 ? E1hpw6[20] : B74iu6);
assign Qyvhu6 = (Qf7iu6 ? E1hpw6[19] : U64iu6);
assign Jyvhu6 = (Qf7iu6 ? E1hpw6[18] : N64iu6);
assign Cyvhu6 = (Qf7iu6 ? E1hpw6[17] : G64iu6);
assign Vxvhu6 = (Qf7iu6 ? E1hpw6[16] : Z54iu6);
assign Oxvhu6 = (Qf7iu6 ? E1hpw6[15] : S54iu6);
assign Hxvhu6 = (Qf7iu6 ? E1hpw6[14] : L54iu6);
assign Axvhu6 = (Qf7iu6 ? E1hpw6[13] : E54iu6);
assign Twvhu6 = (Qf7iu6 ? E1hpw6[12] : X44iu6);
assign Mwvhu6 = (Qf7iu6 ? E1hpw6[11] : Q44iu6);
assign Fwvhu6 = (Qf7iu6 ? E1hpw6[10] : J44iu6);
assign Yvvhu6 = (Qf7iu6 ? E1hpw6[9] : Ym4iu6);
assign Rvvhu6 = (Qf7iu6 ? E1hpw6[8] : Pl4iu6);
assign Kvvhu6 = (Qf7iu6 ? E1hpw6[7] : Gk4iu6);
assign Dvvhu6 = (Qf7iu6 ? E1hpw6[6] : Xi4iu6);
assign Wuvhu6 = (Qf7iu6 ? E1hpw6[5] : Oh4iu6);
assign Puvhu6 = (Qf7iu6 ? E1hpw6[4] : H34iu6);
assign Iuvhu6 = (Qf7iu6 ? E1hpw6[3] : Df4iu6);
assign Buvhu6 = (Qf7iu6 ? E1hpw6[2] : Ud4iu6);
assign Utvhu6 = (Qf7iu6 ? Pzgpw6[1] : O34iu6);
assign Qf7iu6 = (~(A2nhu6 & Zt1iu6));
assign Ntvhu6 = (Xf7iu6 ? R2hpw6[0] : T24iu6);
assign Gtvhu6 = (Xf7iu6 ? R2hpw6[2] : Ud4iu6);
assign Zsvhu6 = (Xf7iu6 ? R2hpw6[1] : O34iu6);
assign Xf7iu6 = (~(Eg7iu6 & A2nhu6));
assign Ssvhu6 = (Lg7iu6 ? G4hpw6[0] : T24iu6);
assign Lsvhu6 = (Lg7iu6 ? G4hpw6[4] : H34iu6);
assign Esvhu6 = (Lg7iu6 ? G4hpw6[3] : Df4iu6);
assign Xrvhu6 = (Lg7iu6 ? G4hpw6[2] : Ud4iu6);
assign Qrvhu6 = (Lg7iu6 ? G4hpw6[1] : O34iu6);
assign Lg7iu6 = (~(Sg7iu6 & A2nhu6));
assign Jrvhu6 = (Zg7iu6 ? V5hpw6[0] : T24iu6);
assign Crvhu6 = (Zg7iu6 ? K7hpw6[31] : Lm1iu6);
assign Vqvhu6 = (Zg7iu6 ? K7hpw6[30] : T94iu6);
assign Oqvhu6 = (Zg7iu6 ? K7hpw6[29] : M94iu6);
assign Hqvhu6 = (Zg7iu6 ? K7hpw6[28] : F94iu6);
assign Aqvhu6 = (Zg7iu6 ? K7hpw6[27] : Y84iu6);
assign Tpvhu6 = (Zg7iu6 ? K7hpw6[26] : R84iu6);
assign Mpvhu6 = (Zg7iu6 ? K7hpw6[25] : K84iu6);
assign Fpvhu6 = (Zg7iu6 ? K7hpw6[24] : D84iu6);
assign Yovhu6 = (Zg7iu6 ? K7hpw6[23] : W74iu6);
assign Rovhu6 = (Zg7iu6 ? K7hpw6[22] : P74iu6);
assign Kovhu6 = (Zg7iu6 ? K7hpw6[21] : I74iu6);
assign Dovhu6 = (Zg7iu6 ? K7hpw6[20] : B74iu6);
assign Wnvhu6 = (Zg7iu6 ? K7hpw6[19] : U64iu6);
assign Pnvhu6 = (Zg7iu6 ? K7hpw6[18] : N64iu6);
assign Invhu6 = (Zg7iu6 ? K7hpw6[17] : G64iu6);
assign Bnvhu6 = (Zg7iu6 ? K7hpw6[16] : Z54iu6);
assign Umvhu6 = (Zg7iu6 ? K7hpw6[15] : S54iu6);
assign Nmvhu6 = (Zg7iu6 ? K7hpw6[14] : L54iu6);
assign Gmvhu6 = (Zg7iu6 ? K7hpw6[13] : E54iu6);
assign Zlvhu6 = (Zg7iu6 ? K7hpw6[12] : X44iu6);
assign Slvhu6 = (Zg7iu6 ? K7hpw6[11] : Q44iu6);
assign Llvhu6 = (Zg7iu6 ? K7hpw6[10] : J44iu6);
assign Elvhu6 = (Zg7iu6 ? K7hpw6[9] : Ym4iu6);
assign Xkvhu6 = (Zg7iu6 ? K7hpw6[8] : Pl4iu6);
assign Qkvhu6 = (Zg7iu6 ? K7hpw6[7] : Gk4iu6);
assign Jkvhu6 = (Zg7iu6 ? K7hpw6[6] : Xi4iu6);
assign Ckvhu6 = (Zg7iu6 ? K7hpw6[5] : Oh4iu6);
assign Vjvhu6 = (Zg7iu6 ? K7hpw6[4] : H34iu6);
assign Ojvhu6 = (Zg7iu6 ? K7hpw6[3] : Df4iu6);
assign Hjvhu6 = (Zg7iu6 ? K7hpw6[2] : Ud4iu6);
assign Ajvhu6 = (Zg7iu6 ? V5hpw6[1] : O34iu6);
assign Zg7iu6 = (~(A2nhu6 & Kw1iu6));
assign Tivhu6 = (~(Gh7iu6 & Nh7iu6));
assign Nh7iu6 = (Uh7iu6 | HREADY);
assign Gh7iu6 = (Bi7iu6 & Ii7iu6);
assign Bi7iu6 = (~(Pi7iu6 & Wi7iu6));
assign Mivhu6 = (Dj7iu6 & Kj7iu6);
assign Kj7iu6 = (Rj7iu6 & Yj7iu6);
assign Rj7iu6 = (~(Xudpw6 & Fk7iu6));
assign Dj7iu6 = (IRQ[0] & Mk7iu6);
assign Mk7iu6 = (~(Tk7iu6 & Al7iu6));
assign Al7iu6 = (Qg6iu6 | Hl7iu6);
assign Fivhu6 = (Ol7iu6 | Vl7iu6);
assign Vl7iu6 = (Ivfhu6 & Cm7iu6);
assign Cm7iu6 = (~(Jm7iu6 & Qm7iu6));
assign Qm7iu6 = (~(Gc5iu6 & Xm7iu6));
assign Xm7iu6 = (Sb5iu6 | Eh6iu6);
assign Yhvhu6 = (En7iu6 | Ln7iu6);
assign En7iu6 = (Zn7iu6 ? Sn7iu6 : Ppfpw6[15]);
assign Sn7iu6 = (HRDATA[15] & Go7iu6);
assign Rhvhu6 = (~(No7iu6 & Uo7iu6));
assign Uo7iu6 = (Bp7iu6 & Ip7iu6);
assign Ip7iu6 = (~(Pp7iu6 & HRDATA[15]));
assign Bp7iu6 = (Wp7iu6 & Dq7iu6);
assign Dq7iu6 = (~(Hrfpw6[15] & Uy4iu6));
assign Wp7iu6 = (~(Kq7iu6 & HRDATA[31]));
assign No7iu6 = (Rq7iu6 & Yq7iu6);
assign Yq7iu6 = (~(Fr7iu6 & Z54iu6));
assign Rq7iu6 = (Mr7iu6 & Tr7iu6);
assign Tr7iu6 = (~(Ppfpw6[15] & A25iu6));
assign Mr7iu6 = (~(R05iu6 & D7fpw6[15]));
assign Khvhu6 = (!As7iu6);
assign As7iu6 = (HREADY ? Os7iu6 : Hs7iu6);
assign Os7iu6 = (~(Vs7iu6 & Ct7iu6));
assign Ct7iu6 = (~(Jt7iu6 & Qt7iu6));
assign Qt7iu6 = (Xt7iu6 & Eu7iu6);
assign Eu7iu6 = (~(Lu7iu6 & Rthhu6));
assign Lu7iu6 = (Smhhu6 & Engpw6[28]);
assign Xt7iu6 = (~(Su7iu6 & Kshhu6));
assign Su7iu6 = (Alhhu6 & Plgpw6[28]);
assign Jt7iu6 = (Zu7iu6 & Gv7iu6);
assign Gv7iu6 = (~(Nv7iu6 & Drhhu6));
assign Nv7iu6 = (Ijhhu6 & Akgpw6[28]);
assign Zu7iu6 = (~(Uv7iu6 & Wphhu6));
assign Uv7iu6 = (Qhhhu6 & Ligpw6[28]);
assign Dhvhu6 = (!Bw7iu6);
assign Bw7iu6 = (HREADY ? Iw7iu6 : Svdpw6);
assign Iw7iu6 = (~(Vs7iu6 & Pw7iu6));
assign Pw7iu6 = (~(Ww7iu6 & Dx7iu6));
assign Dx7iu6 = (Kx7iu6 & Rx7iu6);
assign Rx7iu6 = (~(Yx7iu6 & Rthhu6));
assign Yx7iu6 = (Smhhu6 & Engpw6[27]);
assign Kx7iu6 = (~(Fy7iu6 & Kshhu6));
assign Fy7iu6 = (Alhhu6 & Plgpw6[27]);
assign Ww7iu6 = (My7iu6 & Ty7iu6);
assign Ty7iu6 = (~(Az7iu6 & Drhhu6));
assign Az7iu6 = (Ijhhu6 & Akgpw6[27]);
assign My7iu6 = (~(Hz7iu6 & Wphhu6));
assign Hz7iu6 = (Qhhhu6 & Ligpw6[27]);
assign Vs7iu6 = (Oz7iu6 & Vz7iu6);
assign Vz7iu6 = (~(C08iu6 | Dx0iu6));
assign C08iu6 = (~(Jehhu6 & J08iu6));
assign J08iu6 = (~(Q08iu6 & X08iu6));
assign X08iu6 = (~(E18iu6 & L18iu6));
assign E18iu6 = (S18iu6 & Z18iu6);
assign Oz7iu6 = (~(G28iu6 | Ef1iu6));
assign G28iu6 = (N28iu6 | Rx0iu6);
assign N28iu6 = (!Kohhu6);
assign Wgvhu6 = (~(U28iu6 & B38iu6));
assign B38iu6 = (I38iu6 & P38iu6);
assign P38iu6 = (~(HRDATA[13] & Pp7iu6));
assign I38iu6 = (W38iu6 & D48iu6);
assign D48iu6 = (~(Hrfpw6[13] & Uy4iu6));
assign W38iu6 = (~(HRDATA[29] & Kq7iu6));
assign U28iu6 = (K48iu6 & R48iu6);
assign R48iu6 = (~(A25iu6 & Ppfpw6[13]));
assign K48iu6 = (~(R05iu6 & D7fpw6[13]));
assign Pgvhu6 = (F58iu6 ? S8fpw6[0] : Y48iu6);
assign Y48iu6 = (~(M58iu6 & T58iu6));
assign T58iu6 = (A68iu6 & H68iu6);
assign H68iu6 = (O68iu6 & V68iu6);
assign O68iu6 = (~(C78iu6 | Bi0iu6));
assign A68iu6 = (J78iu6 & Q78iu6);
assign Q78iu6 = (~(X78iu6 & E88iu6));
assign X78iu6 = (L88iu6 ^ S88iu6);
assign J78iu6 = (Z88iu6 & G98iu6);
assign G98iu6 = (~(N98iu6 & U98iu6));
assign N98iu6 = (~(Tr0iu6 | Cyfpw6[6]));
assign Z88iu6 = (~(Ba8iu6 & Ia8iu6));
assign M58iu6 = (Pa8iu6 & Wa8iu6);
assign Wa8iu6 = (Db8iu6 & Kb8iu6);
assign Kb8iu6 = (Rb8iu6 | Yb8iu6);
assign Db8iu6 = (Fc8iu6 & Mc8iu6);
assign Mc8iu6 = (~(Tc8iu6 & Ppfpw6[0]));
assign Fc8iu6 = (Ad8iu6 | Hd8iu6);
assign Pa8iu6 = (Od8iu6 & Vd8iu6);
assign Vd8iu6 = (~(Ce8iu6 & Je8iu6));
assign Od8iu6 = (~(Qe8iu6 & Xe8iu6));
assign Igvhu6 = (Lf8iu6 ? vis_r0_o[4] : Ef8iu6);
assign Bgvhu6 = (Zf8iu6 ? Sf8iu6 : vis_apsr_o[1]);
assign Zf8iu6 = (HREADY & Gg8iu6);
assign Gg8iu6 = (~(Ng8iu6 & Ug8iu6));
assign Sf8iu6 = (~(Bh8iu6 & Ih8iu6));
assign Ih8iu6 = (~(Ph8iu6 & Wh8iu6));
assign Bh8iu6 = (Di8iu6 & Ki8iu6);
assign Ki8iu6 = (~(Ug8iu6 & Ri8iu6));
assign Di8iu6 = (~(Yi8iu6 & Fj8iu6));
assign Ufvhu6 = (~(Mj8iu6 & Tj8iu6));
assign Tj8iu6 = (Ak8iu6 & Hk8iu6);
assign Hk8iu6 = (~(Ok8iu6 & vis_pc_o[28]));
assign Ak8iu6 = (Vk8iu6 & Cl8iu6);
assign Cl8iu6 = (~(Jl8iu6 & Dx0iu6));
assign Vk8iu6 = (~(Ql8iu6 & vis_apsr_o[1]));
assign Mj8iu6 = (Xl8iu6 & Em8iu6);
assign Em8iu6 = (Lm8iu6 | Sm8iu6);
assign Xl8iu6 = (~(Zm8iu6 & M94iu6));
assign Nfvhu6 = (Nn8iu6 ? vis_tbit_o : Gn8iu6);
assign Nn8iu6 = (Un8iu6 & Bo8iu6);
assign Bo8iu6 = (~(Io8iu6 & Po8iu6));
assign Po8iu6 = (Wo8iu6 & Dp8iu6);
assign Wo8iu6 = (~(Kp8iu6 & Rp8iu6));
assign Rp8iu6 = (~(Yp8iu6 | Fq8iu6));
assign Kp8iu6 = (Mq8iu6 & Tq8iu6);
assign Tq8iu6 = (Mr0iu6 | Tr0iu6);
assign Mq8iu6 = (Cyfpw6[3] | Y7ghu6);
assign Io8iu6 = (Ar8iu6 & Hr8iu6);
assign Un8iu6 = (~(HREADY & Or8iu6));
assign Or8iu6 = (~(Vr8iu6 & Cs8iu6));
assign Gn8iu6 = (Vr8iu6 ? Js8iu6 : Fkfpw6[24]);
assign Js8iu6 = (~(Qs8iu6 & Xs8iu6));
assign Xs8iu6 = (~(Eafpw6[0] & Et8iu6));
assign Qs8iu6 = (Lt8iu6 & St8iu6);
assign St8iu6 = (Zt8iu6 | Gu8iu6);
assign Lt8iu6 = (~(Yi8iu6 & Nu8iu6));
assign Gfvhu6 = (~(Uu8iu6 & Bv8iu6));
assign Bv8iu6 = (Iv8iu6 & Pv8iu6);
assign Pv8iu6 = (~(Hrfpw6[14] & Uy4iu6));
assign Iv8iu6 = (Wv8iu6 & Dw8iu6);
assign Dw8iu6 = (~(M15iu6 & Kw8iu6));
assign Wv8iu6 = (~(Pz4iu6 & Rw8iu6));
assign Uu8iu6 = (Yw8iu6 & Fx8iu6);
assign Fx8iu6 = (~(Ppfpw6[14] & A25iu6));
assign Yw8iu6 = (~(R05iu6 & D7fpw6[14]));
assign Zevhu6 = (Mx8iu6 ? vis_r1_o[4] : Ef8iu6);
assign Sevhu6 = (Mx8iu6 ? vis_r1_o[0] : Tx8iu6);
assign Levhu6 = (Hy8iu6 ? Ay8iu6 : Iwfpw6[0]);
assign Eevhu6 = (Lf8iu6 ? vis_r0_o[0] : Tx8iu6);
assign Xdvhu6 = (Vy8iu6 ? Oy8iu6 : vis_primask_o);
assign Vy8iu6 = (~(Eh6iu6 | Cz8iu6));
assign Qdvhu6 = (~(Jz8iu6 & Qz8iu6));
assign Qz8iu6 = (Xz8iu6 & E09iu6);
assign E09iu6 = (~(Ql8iu6 & vis_ipsr_o[0]));
assign Xz8iu6 = (L09iu6 & S09iu6);
assign S09iu6 = (~(Jl8iu6 & Z09iu6));
assign Z09iu6 = (Ay8iu6 | G19iu6);
assign G19iu6 = (~(N19iu6 | U19iu6));
assign L09iu6 = (~(B29iu6 & vis_primask_o));
assign Jz8iu6 = (I29iu6 & P29iu6);
assign P29iu6 = (~(W29iu6 & Fkfpw6[0]));
assign I29iu6 = (~(Zm8iu6 & T24iu6));
assign Jdvhu6 = (Mx8iu6 ? vis_r1_o[31] : D39iu6);
assign Cdvhu6 = (Lf8iu6 ? vis_r0_o[31] : D39iu6);
assign Vcvhu6 = (Mx8iu6 ? vis_r1_o[30] : K39iu6);
assign Ocvhu6 = (Lf8iu6 ? vis_r0_o[30] : K39iu6);
assign Hcvhu6 = (~(R39iu6 & Y39iu6));
assign Y39iu6 = (~(Jfgpw6[1] & Eh6iu6));
assign R39iu6 = (F49iu6 & Ii7iu6);
assign F49iu6 = (~(M49iu6 & Wi7iu6));
assign Acvhu6 = (~(T49iu6 & A59iu6));
assign A59iu6 = (~(Vbgpw6[31] & H59iu6));
assign H59iu6 = (~(HWDATA[31] & O59iu6));
assign T49iu6 = (~(V59iu6 & HWDATA[31]));
assign Tbvhu6 = (~(C69iu6 & J69iu6));
assign J69iu6 = (~(Vbgpw6[0] & Q69iu6));
assign Q69iu6 = (~(HWDATA[0] & O59iu6));
assign C69iu6 = (~(V59iu6 & HWDATA[0]));
assign Mbvhu6 = (~(X69iu6 & E79iu6));
assign E79iu6 = (~(Jfgpw6[3] & Eh6iu6));
assign X69iu6 = (L79iu6 & Ii7iu6);
assign L79iu6 = (~(S79iu6 & Wi7iu6));
assign S79iu6 = (~(HADDR[3] ^ Z79iu6));
assign Fbvhu6 = (~(G89iu6 & N89iu6));
assign N89iu6 = (U89iu6 | HREADY);
assign G89iu6 = (B99iu6 & Ii7iu6);
assign B99iu6 = (~(I99iu6 & Wi7iu6));
assign I99iu6 = (~(HADDR[2] ^ P99iu6));
assign Yavhu6 = (~(W99iu6 & Da9iu6));
assign Da9iu6 = (Ka9iu6 | HREADY);
assign W99iu6 = (Ra9iu6 & Ii7iu6);
assign Ii7iu6 = (~(Wi7iu6 & Ya9iu6));
assign Ya9iu6 = (~(Fb9iu6 & Mb9iu6));
assign Mb9iu6 = (HSIZE[1] & Tb9iu6);
assign Tb9iu6 = (~(Ac9iu6 & Hc9iu6));
assign Hc9iu6 = (~(Oc9iu6 & Vc9iu6));
assign Vc9iu6 = (~(Cd9iu6 | HADDR[9]));
assign Cd9iu6 = (~(Jd9iu6 & Qd9iu6));
assign Qd9iu6 = (~(HADDR[6] & Xd9iu6));
assign Xd9iu6 = (~(HADDR[7] & Ee9iu6));
assign Ee9iu6 = (HADDR[3] | HADDR[2]);
assign Jd9iu6 = (~(HADDR[7] & Le9iu6));
assign Le9iu6 = (~(Se9iu6 & HADDR[11]));
assign Se9iu6 = (~(M49iu6 | Ze9iu6));
assign Oc9iu6 = (Gf9iu6 & Nf9iu6);
assign Nf9iu6 = (HADDR[11] ? Uf9iu6 : Pi7iu6);
assign Uf9iu6 = (Bg9iu6 & Ig9iu6);
assign Ig9iu6 = (Pg9iu6 & Wg9iu6);
assign Wg9iu6 = (~(HADDR[3] & Dh9iu6));
assign Dh9iu6 = (M49iu6 | HADDR[2]);
assign Pg9iu6 = (M49iu6 | HADDR[6]);
assign M49iu6 = (!HADDR[4]);
assign Bg9iu6 = (HADDR[5] & Kh9iu6);
assign Kh9iu6 = (Rh9iu6 | Xg6iu6);
assign Rh9iu6 = (!HADDR[2]);
assign Gf9iu6 = (HADDR[10] & Yh9iu6);
assign Yh9iu6 = (Z79iu6 | HADDR[8]);
assign Ac9iu6 = (HADDR[11] ? Mi9iu6 : Fi9iu6);
assign HADDR[11] = (Ze9iu6 ? Tugpw6[9] : Jshpw6[11]);
assign Mi9iu6 = (~(Ti9iu6 & Aj9iu6));
assign Aj9iu6 = (Hj9iu6 & Oj9iu6);
assign Oj9iu6 = (HADDR[10] & Vj9iu6);
assign Vj9iu6 = (Ck9iu6 | HADDR[2]);
assign Hj9iu6 = (~(HADDR[6] | Pi7iu6));
assign Ti9iu6 = (Jk9iu6 & P99iu6);
assign P99iu6 = (!HADDR[7]);
assign Jk9iu6 = (~(HADDR[9] | HADDR[5]));
assign Fi9iu6 = (~(Qk9iu6 & Z79iu6));
assign Z79iu6 = (!HADDR[5]);
assign HADDR[5] = (Xg6iu6 ? Jshpw6[5] : Tugpw6[3]);
assign Qk9iu6 = (Xk9iu6 & El9iu6);
assign El9iu6 = (!HADDR[6]);
assign Xk9iu6 = (Zl9iu6 ? Sl9iu6 : Ll9iu6);
assign Zl9iu6 = (~(HADDR[4] | HADDR[3]));
assign HADDR[4] = (Xg6iu6 ? Jshpw6[4] : Tugpw6[2]);
assign Sl9iu6 = (Gm9iu6 & Nm9iu6);
assign Nm9iu6 = (~(HADDR[9] ^ Pi7iu6));
assign Gm9iu6 = (~(HADDR[2] | HADDR[10]));
assign HADDR[2] = (Xg6iu6 ? P47iu6 : Tugpw6[0]);
assign P47iu6 = (Wqzhu6 ? Vo4iu6 : Tnhpw6[2]);
assign Ll9iu6 = (Um9iu6 & Pi7iu6);
assign Pi7iu6 = (!HADDR[8]);
assign HADDR[8] = (Xg6iu6 ? Jshpw6[8] : Tugpw6[6]);
assign Um9iu6 = (~(HADDR[9] | HADDR[7]));
assign HADDR[7] = (Xg6iu6 ? Jshpw6[7] : Tugpw6[5]);
assign Fb9iu6 = (Bn9iu6 & HADDR[15]);
assign Bn9iu6 = (Xg6iu6 ? Pn9iu6 : In9iu6);
assign Pn9iu6 = (Wn9iu6 & Fs6iu6);
assign Fs6iu6 = (Do9iu6 & Ko9iu6);
assign Ko9iu6 = (Ro9iu6 & Yo9iu6);
assign Yo9iu6 = (!Jshpw6[25]);
assign Ro9iu6 = (~(Jshpw6[26] | Jshpw6[27]));
assign Do9iu6 = (Fp9iu6 & Mp9iu6);
assign Mp9iu6 = (!Jshpw6[22]);
assign Fp9iu6 = (~(Jshpw6[23] | Jshpw6[24]));
assign Wn9iu6 = (Tp9iu6 & Aq9iu6);
assign Aq9iu6 = (At6iu6 & Bx6iu6);
assign Bx6iu6 = (!Jshpw6[12]);
assign At6iu6 = (~(Jshpw6[20] | Jshpw6[21]));
assign Tp9iu6 = (Kc7iu6 & Mz6iu6);
assign Mz6iu6 = (Hq9iu6 & Oq9iu6);
assign Oq9iu6 = (~(Jshpw6[18] | Jshpw6[19]));
assign Hq9iu6 = (~(Jshpw6[16] | Jshpw6[17]));
assign Kc7iu6 = (Jshpw6[14] & Jshpw6[13]);
assign In9iu6 = (Vq9iu6 & Cr9iu6);
assign Cr9iu6 = (Jr9iu6 & Qr9iu6);
assign Qr9iu6 = (Xr9iu6 & Es9iu6);
assign Es9iu6 = (~(Pxdpw6 | Ixdpw6));
assign Xr9iu6 = (~(Dydpw6 | Wxdpw6));
assign Jr9iu6 = (Ls9iu6 & Ss9iu6);
assign Ss9iu6 = (~(Rydpw6 | Kydpw6));
assign Ls9iu6 = (~(Fzdpw6 | Yydpw6));
assign Vq9iu6 = (Zs9iu6 & Gt9iu6);
assign Gt9iu6 = (Nt9iu6 & Ut9iu6);
assign Ut9iu6 = (~(Tzdpw6 | Mzdpw6));
assign Nt9iu6 = (~(H0epw6 | A0epw6));
assign Zs9iu6 = (Bu9iu6 & Tugpw6[12]);
assign Bu9iu6 = (~(Iu9iu6 | O0epw6));
assign Iu9iu6 = (!Tugpw6[11]);
assign Ra9iu6 = (~(Pu9iu6 & Wi7iu6));
assign Pu9iu6 = (~(HADDR[10] ^ Ck9iu6));
assign Ck9iu6 = (!HADDR[3]);
assign HADDR[3] = (Xg6iu6 ? I47iu6 : Tugpw6[1]);
assign I47iu6 = (Wqzhu6 ? Wu9iu6 : Tnhpw6[3]);
assign HADDR[10] = (Xg6iu6 ? Jshpw6[10] : Tugpw6[8]);
assign Ravhu6 = (Dv9iu6 ? R4gpw6[7] : HWDATA[31]);
assign Kavhu6 = (~(Kv9iu6 & Rv9iu6));
assign Rv9iu6 = (Yv9iu6 & Fw9iu6);
assign Fw9iu6 = (~(Jl8iu6 & Mzdpw6));
assign Yv9iu6 = (~(vis_pc_o[22] & Ok8iu6));
assign Kv9iu6 = (Mw9iu6 & Tw9iu6);
assign Tw9iu6 = (Lm8iu6 | Ax9iu6);
assign Mw9iu6 = (Hx9iu6 | Ox9iu6);
assign Davhu6 = (Mx8iu6 ? vis_r1_o[23] : Vx9iu6);
assign W9vhu6 = (Lf8iu6 ? vis_r0_o[23] : Vx9iu6);
assign P9vhu6 = (Jy9iu6 ? Cy9iu6 : Vrfhu6);
assign Jy9iu6 = (HREADY & Qy9iu6);
assign Qy9iu6 = (~(Xy9iu6 & Ez9iu6));
assign Ez9iu6 = (Lz9iu6 & Sz9iu6);
assign Sz9iu6 = (Zz9iu6 & G0aiu6);
assign G0aiu6 = (~(N0aiu6 & U0aiu6));
assign N0aiu6 = (~(Cyfpw6[6] | Y7ghu6));
assign Zz9iu6 = (B1aiu6 & I1aiu6);
assign Lz9iu6 = (P1aiu6 & W1aiu6);
assign W1aiu6 = (~(D2aiu6 & K2aiu6));
assign D2aiu6 = (~(R2aiu6 | Cyfpw6[4]));
assign P1aiu6 = (~(Y2aiu6 & F3aiu6));
assign Xy9iu6 = (M3aiu6 & T3aiu6);
assign T3aiu6 = (A4aiu6 & H4aiu6);
assign H4aiu6 = (O4aiu6 | V4aiu6);
assign A4aiu6 = (C5aiu6 & J5aiu6);
assign C5aiu6 = (Q5aiu6 | X5aiu6);
assign M3aiu6 = (E6aiu6 & L6aiu6);
assign E6aiu6 = (~(S6aiu6 & Z6aiu6));
assign Cy9iu6 = (~(G7aiu6 & N7aiu6));
assign N7aiu6 = (~(U7aiu6 & B8aiu6));
assign B8aiu6 = (I8aiu6 | P8aiu6);
assign P8aiu6 = (Cyfpw6[3] ? D9aiu6 : W8aiu6);
assign D9aiu6 = (K9aiu6 | R9aiu6);
assign I8aiu6 = (~(Y9aiu6 & Faaiu6));
assign Y9aiu6 = (Mr0iu6 ? D7fpw6[3] : Cyfpw6[5]);
assign U7aiu6 = (vis_control_o | Maaiu6);
assign Maaiu6 = (~(Taaiu6 | Quzhu6));
assign G7aiu6 = (Cyfpw6[3] ? Hbaiu6 : Abaiu6);
assign Hbaiu6 = (~(Obaiu6 & Vbaiu6));
assign Vbaiu6 = (~(R2aiu6 | D7fpw6[0]));
assign Obaiu6 = (~(Ccaiu6 | V4aiu6));
assign Abaiu6 = (Rb8iu6 | Jcaiu6);
assign I9vhu6 = (Mx8iu6 ? vis_r1_o[2] : Qcaiu6);
assign B9vhu6 = (Lf8iu6 ? vis_r0_o[2] : Qcaiu6);
assign U8vhu6 = (~(Xcaiu6 & Edaiu6));
assign Edaiu6 = (~(Ldaiu6 & Hy8iu6));
assign Ldaiu6 = (~(Z18iu6 | Sdaiu6));
assign Xcaiu6 = (~(Zdaiu6 & Eh6iu6));
assign Zdaiu6 = (~(Geaiu6 & Neaiu6));
assign Neaiu6 = (~(V3xhu6 & Ueaiu6));
assign Ueaiu6 = (~(Bfaiu6 & Ifaiu6));
assign Ifaiu6 = (Pfaiu6 & Wfaiu6);
assign Wfaiu6 = (~(K2aiu6 & Dgaiu6));
assign Dgaiu6 = (~(Kgaiu6 & Rgaiu6));
assign Rgaiu6 = (~(Ygaiu6 & Fhaiu6));
assign Ygaiu6 = (~(As0iu6 | Y7ghu6));
assign Pfaiu6 = (Mhaiu6 & Thaiu6);
assign Mhaiu6 = (~(Aiaiu6 & Hiaiu6));
assign Aiaiu6 = (Oiaiu6 & Viaiu6);
assign Viaiu6 = (~(Cjaiu6 & Jjaiu6));
assign Jjaiu6 = (Qjaiu6 | Cyfpw6[3]);
assign Cjaiu6 = (Xjaiu6 & Ekaiu6);
assign Xjaiu6 = (As0iu6 | Lkaiu6);
assign Bfaiu6 = (Skaiu6 & Zkaiu6);
assign Zkaiu6 = (~(Glaiu6 & Nlaiu6));
assign Skaiu6 = (Ulaiu6 & Bmaiu6);
assign Bmaiu6 = (~(Imaiu6 & Pmaiu6));
assign Pmaiu6 = (~(Wmaiu6 & Dnaiu6));
assign Dnaiu6 = (Knaiu6 | Cyfpw6[1]);
assign Ulaiu6 = (~(Cyfpw6[7] & Rnaiu6));
assign Rnaiu6 = (~(Ynaiu6 & Foaiu6));
assign Foaiu6 = (~(Moaiu6 & Ii0iu6));
assign Ynaiu6 = (~(Toaiu6 & Apaiu6));
assign N8vhu6 = (~(Hpaiu6 & Opaiu6));
assign Opaiu6 = (~(Vpaiu6 & Cqaiu6));
assign Vpaiu6 = (~(Jqaiu6 & Qqaiu6));
assign Qqaiu6 = (Xqaiu6 & Eraiu6);
assign Eraiu6 = (~(Lraiu6 & Ja5iu6));
assign Xqaiu6 = (Sraiu6 & Zraiu6);
assign Sraiu6 = (~(Gsaiu6 & Nsaiu6));
assign Jqaiu6 = (Usaiu6 & HREADY);
assign Hpaiu6 = (~(SLEEPHOLDREQn & HREADY));
assign G8vhu6 = (~(Li5iu6 & Btaiu6));
assign Btaiu6 = (~(Itaiu6 & Righu6));
assign Itaiu6 = (~(Ptaiu6 | Qg6iu6));
assign Li5iu6 = (Wtaiu6 & Duaiu6);
assign Duaiu6 = (~(Kuaiu6 & Ruaiu6));
assign Kuaiu6 = (~(Yuaiu6 & Fvaiu6));
assign Fvaiu6 = (Mvaiu6 & Tvaiu6);
assign Tvaiu6 = (~(Awaiu6 & Hwaiu6));
assign Awaiu6 = (~(Owaiu6 | Vwaiu6));
assign Mvaiu6 = (~(Cxaiu6 & Jxaiu6));
assign Cxaiu6 = (~(Qxaiu6 | D7fpw6[14]));
assign Yuaiu6 = (Xxaiu6 & Eyaiu6);
assign Eyaiu6 = (~(Lyaiu6 & L3ehu6));
assign Wtaiu6 = (Syaiu6 & Zyaiu6);
assign Zyaiu6 = (~(Lyaiu6 & Gzaiu6));
assign Gzaiu6 = (~(Nzaiu6 | L3ehu6));
assign Nzaiu6 = (Uzaiu6 & B0biu6);
assign Lyaiu6 = (~(K9aiu6 | Geaiu6));
assign Syaiu6 = (I0biu6 | P0biu6);
assign Z7vhu6 = (~(W0biu6 & D1biu6));
assign D1biu6 = (~(K1biu6 & R1biu6));
assign R1biu6 = (~(Geaiu6 | L3ehu6));
assign K1biu6 = (Y1biu6 & F2biu6);
assign Y1biu6 = (Uzaiu6 ? M2biu6 : Quzhu6);
assign W0biu6 = (~(Qwdhu6 & T2biu6));
assign S7vhu6 = (~(A3biu6 & H3biu6));
assign H3biu6 = (O3biu6 & V3biu6);
assign V3biu6 = (~(HRDATA[0] & Pp7iu6));
assign O3biu6 = (C4biu6 & J4biu6);
assign J4biu6 = (~(Hrfpw6[0] & Uy4iu6));
assign C4biu6 = (~(HRDATA[16] & Kq7iu6));
assign A3biu6 = (Q4biu6 & X4biu6);
assign X4biu6 = (~(Fr7iu6 & T24iu6));
assign Q4biu6 = (E5biu6 & L5biu6);
assign L5biu6 = (~(Ppfpw6[0] & A25iu6));
assign E5biu6 = (~(R05iu6 & D7fpw6[0]));
assign L7vhu6 = (F58iu6 ? S8fpw6[1] : S5biu6);
assign S5biu6 = (~(Z5biu6 & G6biu6));
assign G6biu6 = (N6biu6 & U6biu6);
assign U6biu6 = (B7biu6 & V68iu6);
assign B7biu6 = (~(I7biu6 & E88iu6));
assign I7biu6 = (P7biu6 ^ W7biu6);
assign N6biu6 = (D8biu6 & K8biu6);
assign K8biu6 = (~(R8biu6 & Ce8iu6));
assign R8biu6 = (~(Y8biu6 ^ S8fpw6[0]));
assign D8biu6 = (~(Tc8iu6 & Ppfpw6[1]));
assign Z5biu6 = (F9biu6 & M9biu6);
assign M9biu6 = (T9biu6 & Aabiu6);
assign Aabiu6 = (O95iu6 | Hd8iu6);
assign T9biu6 = (~(Habiu6 & D7fpw6[0]));
assign F9biu6 = (Oabiu6 & Vabiu6);
assign Vabiu6 = (Ccaiu6 | Yb8iu6);
assign Oabiu6 = (~(Cbbiu6 & D7fpw6[6]));
assign E7vhu6 = (~(Jbbiu6 & Qbbiu6));
assign Qbbiu6 = (~(D8hhu6 & Xbbiu6));
assign X6vhu6 = (~(Qw4iu6 & Ecbiu6));
assign Ecbiu6 = (~(Dhgpw6[1] & Lcbiu6));
assign Lcbiu6 = (~(Scbiu6 & O34iu6));
assign Qw4iu6 = (~(W8aiu6 & Cyfpw6[0]));
assign Q6vhu6 = (Zcbiu6 & Gdbiu6);
assign Gdbiu6 = (Ndbiu6 & Udbiu6);
assign Ndbiu6 = (~(Npdpw6 & Bebiu6));
assign Zcbiu6 = (IRQ[31] & Iebiu6);
assign Iebiu6 = (~(Tk7iu6 & Pebiu6));
assign Pebiu6 = (Webiu6 | Qg6iu6);
assign J6vhu6 = (Dfbiu6 & Kfbiu6);
assign Kfbiu6 = (Rfbiu6 & Yfbiu6);
assign Rfbiu6 = (~(Updpw6 & Fgbiu6));
assign Dfbiu6 = (IRQ[29] & Mgbiu6);
assign Mgbiu6 = (~(Tk7iu6 & Tgbiu6));
assign Tgbiu6 = (Qg6iu6 | Ahbiu6);
assign C6vhu6 = (~(Hhbiu6 & Ohbiu6));
assign Ohbiu6 = (Vhbiu6 | Cibiu6);
assign Hhbiu6 = (Jibiu6 & Qibiu6);
assign Qibiu6 = (~(Xibiu6 & Ppfpw6[5]));
assign Jibiu6 = (Ejbiu6 | Ljbiu6);
assign V5vhu6 = (~(Sjbiu6 & Zjbiu6));
assign Zjbiu6 = (Gkbiu6 & Nkbiu6);
assign Nkbiu6 = (~(HRDATA[8] & Pp7iu6));
assign Gkbiu6 = (Ukbiu6 & Blbiu6);
assign Blbiu6 = (~(Hrfpw6[8] & Uy4iu6));
assign Ukbiu6 = (~(HRDATA[24] & Kq7iu6));
assign Sjbiu6 = (Ilbiu6 & Plbiu6);
assign Plbiu6 = (~(A25iu6 & Ppfpw6[8]));
assign Ilbiu6 = (~(D7fpw6[8] & R05iu6));
assign O5vhu6 = (~(Wlbiu6 & Dmbiu6));
assign Dmbiu6 = (Jm7iu6 | Kmbiu6);
assign Wlbiu6 = (Rmbiu6 & Ymbiu6);
assign Ymbiu6 = (~(Ppfpw6[0] & Fnbiu6));
assign Rmbiu6 = (~(Mnbiu6 & HRDATA[0]));
assign H5vhu6 = (~(Tnbiu6 & Aobiu6));
assign Aobiu6 = (~(Hobiu6 & Kw8iu6));
assign Kw8iu6 = (~(Svdpw6 & Oobiu6));
assign Oobiu6 = (~(HRDATA[14] & Vobiu6));
assign Tnbiu6 = (~(Ppfpw6[14] & Cpbiu6));
assign A5vhu6 = (~(Jpbiu6 & Qpbiu6));
assign Qpbiu6 = (Xpbiu6 & Eqbiu6);
assign Eqbiu6 = (~(Xlfpw6[8] & Lqbiu6));
assign Xpbiu6 = (~(IRQLATENCY[7] & Ol7iu6));
assign Jpbiu6 = (Sqbiu6 & Zqbiu6);
assign Zqbiu6 = (~(Mnbiu6 & HRDATA[13]));
assign Sqbiu6 = (~(Cpbiu6 & Ppfpw6[13]));
assign T4vhu6 = (~(Grbiu6 & Nrbiu6));
assign Nrbiu6 = (Urbiu6 & Bsbiu6);
assign Bsbiu6 = (~(Xlfpw6[7] & Lqbiu6));
assign Urbiu6 = (~(IRQLATENCY[6] & Ol7iu6));
assign Grbiu6 = (Isbiu6 & Psbiu6);
assign Psbiu6 = (~(Mnbiu6 & HRDATA[12]));
assign Isbiu6 = (~(Cpbiu6 & Ppfpw6[12]));
assign M4vhu6 = (~(Wsbiu6 & Dtbiu6));
assign Dtbiu6 = (Ktbiu6 & Rtbiu6);
assign Rtbiu6 = (~(Xlfpw6[6] & Lqbiu6));
assign Ktbiu6 = (~(IRQLATENCY[5] & Ol7iu6));
assign Wsbiu6 = (Ytbiu6 & Fubiu6);
assign Fubiu6 = (~(HRDATA[11] & Mnbiu6));
assign Ytbiu6 = (~(Cpbiu6 & Ppfpw6[11]));
assign F4vhu6 = (~(Mubiu6 & Tubiu6));
assign Tubiu6 = (Avbiu6 & Hvbiu6);
assign Hvbiu6 = (~(Xlfpw6[5] & Lqbiu6));
assign Avbiu6 = (~(IRQLATENCY[4] & Ol7iu6));
assign Mubiu6 = (Ovbiu6 & Vvbiu6);
assign Vvbiu6 = (~(Mnbiu6 & HRDATA[10]));
assign Ovbiu6 = (~(Cpbiu6 & Ppfpw6[10]));
assign Y3vhu6 = (~(Cwbiu6 & Jwbiu6));
assign Jwbiu6 = (Qwbiu6 & Xwbiu6);
assign Xwbiu6 = (~(Xlfpw6[4] & Lqbiu6));
assign Qwbiu6 = (~(IRQLATENCY[3] & Ol7iu6));
assign Cwbiu6 = (Exbiu6 & Lxbiu6);
assign Lxbiu6 = (~(HRDATA[9] & Mnbiu6));
assign Exbiu6 = (~(Cpbiu6 & Ppfpw6[9]));
assign R3vhu6 = (~(Sxbiu6 & Zxbiu6));
assign Zxbiu6 = (Gybiu6 & Nybiu6);
assign Nybiu6 = (~(Xlfpw6[3] & Lqbiu6));
assign Gybiu6 = (~(IRQLATENCY[2] & Ol7iu6));
assign Sxbiu6 = (Uybiu6 & Bzbiu6);
assign Bzbiu6 = (~(Mnbiu6 & HRDATA[8]));
assign Uybiu6 = (~(Cpbiu6 & Ppfpw6[8]));
assign K3vhu6 = (~(Izbiu6 & Pzbiu6));
assign Pzbiu6 = (Wzbiu6 & D0ciu6);
assign D0ciu6 = (~(Xlfpw6[2] & Lqbiu6));
assign Wzbiu6 = (~(IRQLATENCY[1] & Ol7iu6));
assign Izbiu6 = (K0ciu6 & R0ciu6);
assign R0ciu6 = (~(Mnbiu6 & HRDATA[7]));
assign K0ciu6 = (~(Cpbiu6 & Ppfpw6[7]));
assign D3vhu6 = (~(Y0ciu6 & F1ciu6));
assign F1ciu6 = (M1ciu6 & T1ciu6);
assign T1ciu6 = (~(Xlfpw6[1] & Lqbiu6));
assign Lqbiu6 = (~(Ol7iu6 | A2ciu6));
assign M1ciu6 = (~(IRQLATENCY[0] & Ol7iu6));
assign Ol7iu6 = (H2ciu6 & O2ciu6);
assign O2ciu6 = (~(V2ciu6 & C3ciu6));
assign C3ciu6 = (J3ciu6 & Q3ciu6);
assign Q3ciu6 = (Ivfhu6 & X3ciu6);
assign X3ciu6 = (~(Ppfpw6[1] ^ E4ciu6));
assign J3ciu6 = (L4ciu6 & S4ciu6);
assign S4ciu6 = (Z4ciu6 ^ Ppfpw6[4]);
assign L4ciu6 = (Kmbiu6 ^ Ppfpw6[0]);
assign V2ciu6 = (G5ciu6 & N5ciu6);
assign N5ciu6 = (U5ciu6 ^ Ppfpw6[2]);
assign G5ciu6 = (B6ciu6 & I6ciu6);
assign I6ciu6 = (P6ciu6 ^ Ppfpw6[3]);
assign B6ciu6 = (W6ciu6 ^ Ppfpw6[5]);
assign Y0ciu6 = (D7ciu6 & K7ciu6);
assign K7ciu6 = (~(Mnbiu6 & HRDATA[6]));
assign D7ciu6 = (~(Cpbiu6 & Ppfpw6[6]));
assign W2vhu6 = (~(R7ciu6 & Y7ciu6));
assign Y7ciu6 = (~(vis_ipsr_o[0] & F8ciu6));
assign R7ciu6 = (M8ciu6 & T8ciu6);
assign T8ciu6 = (~(Xibiu6 & Ppfpw6[0]));
assign M8ciu6 = (Ejbiu6 | Zt8iu6);
assign P2vhu6 = (~(A9ciu6 & H9ciu6));
assign H9ciu6 = (~(O9ciu6 & H2ciu6));
assign O9ciu6 = (HREADY & V9ciu6);
assign A9ciu6 = (~(Fvdhu6 & Caciu6));
assign Caciu6 = (~(HREADY & Jaciu6));
assign Jaciu6 = (~(Gc5iu6 & V9ciu6));
assign V9ciu6 = (Uzaiu6 | Qaciu6);
assign I2vhu6 = (~(Xaciu6 & Ebciu6));
assign Ebciu6 = (Jm7iu6 | W6ciu6);
assign Xaciu6 = (Lbciu6 & Sbciu6);
assign Sbciu6 = (~(Ppfpw6[5] & Fnbiu6));
assign Lbciu6 = (~(Mnbiu6 & HRDATA[5]));
assign B2vhu6 = (~(Zbciu6 & Gcciu6));
assign Gcciu6 = (Jm7iu6 | Z4ciu6);
assign Zbciu6 = (Ncciu6 & Ucciu6);
assign Ucciu6 = (~(Ppfpw6[4] & Fnbiu6));
assign Ncciu6 = (~(Mnbiu6 & HRDATA[4]));
assign U1vhu6 = (~(Bdciu6 & Idciu6));
assign Idciu6 = (Jm7iu6 | P6ciu6);
assign Bdciu6 = (Pdciu6 & Wdciu6);
assign Wdciu6 = (~(Ppfpw6[3] & Fnbiu6));
assign Pdciu6 = (~(HRDATA[3] & Mnbiu6));
assign N1vhu6 = (~(Deciu6 & Keciu6));
assign Keciu6 = (Jm7iu6 | U5ciu6);
assign Deciu6 = (Reciu6 & Yeciu6);
assign Yeciu6 = (~(Ppfpw6[2] & Fnbiu6));
assign Reciu6 = (~(Mnbiu6 & HRDATA[2]));
assign G1vhu6 = (~(Ffciu6 & Mfciu6));
assign Mfciu6 = (Tfciu6 | Cibiu6);
assign Ffciu6 = (Agciu6 & Hgciu6);
assign Hgciu6 = (~(Xibiu6 & Ppfpw6[2]));
assign Agciu6 = (Ejbiu6 | Ogciu6);
assign Z0vhu6 = (~(Vgciu6 & Chciu6));
assign Chciu6 = (~(H2ciu6 & E4ciu6));
assign Vgciu6 = (Jhciu6 & Qhciu6);
assign Qhciu6 = (~(Ppfpw6[1] & Fnbiu6));
assign Fnbiu6 = (~(Zn7iu6 & Xhciu6));
assign Xhciu6 = (A2ciu6 | H2ciu6);
assign Jhciu6 = (~(HRDATA[1] & Mnbiu6));
assign Mnbiu6 = (Hobiu6 & Go7iu6);
assign S0vhu6 = (~(Eiciu6 & Liciu6));
assign Liciu6 = (Siciu6 | Cibiu6);
assign Eiciu6 = (Ziciu6 & Gjciu6);
assign Gjciu6 = (~(Xibiu6 & Ppfpw6[1]));
assign Ziciu6 = (Ejbiu6 | Njciu6);
assign L0vhu6 = (Hobiu6 | Ujciu6);
assign Ujciu6 = (Bkciu6 & Ikciu6);
assign Ikciu6 = (Ntfhu6 & Pkciu6);
assign Bkciu6 = (Cpbiu6 & R05iu6);
assign Hobiu6 = (~(Ln7iu6 | Cpbiu6));
assign Cpbiu6 = (!Zn7iu6);
assign E0vhu6 = (~(Wkciu6 & Dlciu6));
assign Dlciu6 = (Klciu6 & Rlciu6);
assign Rlciu6 = (~(HRDATA[12] & Pp7iu6));
assign Klciu6 = (Ylciu6 & Fmciu6);
assign Fmciu6 = (~(Hrfpw6[12] & Uy4iu6));
assign Ylciu6 = (~(HRDATA[28] & Kq7iu6));
assign Wkciu6 = (Mmciu6 & Tmciu6);
assign Tmciu6 = (~(A25iu6 & Ppfpw6[12]));
assign Mmciu6 = (~(R05iu6 & D7fpw6[12]));
assign Xzuhu6 = (~(Anciu6 & Hnciu6));
assign Hnciu6 = (Onciu6 & Vnciu6);
assign Vnciu6 = (~(HRDATA[11] & Pp7iu6));
assign Onciu6 = (Cociu6 & Jociu6);
assign Jociu6 = (~(Hrfpw6[11] & Uy4iu6));
assign Cociu6 = (~(HRDATA[27] & Kq7iu6));
assign Anciu6 = (Qociu6 & Xociu6);
assign Xociu6 = (~(A25iu6 & Ppfpw6[11]));
assign Qociu6 = (~(R05iu6 & D7fpw6[11]));
assign Qzuhu6 = (~(Epciu6 & Lpciu6));
assign Lpciu6 = (Spciu6 & Zpciu6);
assign Zpciu6 = (~(HRDATA[10] & Pp7iu6));
assign Spciu6 = (Gqciu6 & Nqciu6);
assign Nqciu6 = (~(Hrfpw6[10] & Uy4iu6));
assign Gqciu6 = (~(HRDATA[26] & Kq7iu6));
assign Epciu6 = (Uqciu6 & Brciu6);
assign Brciu6 = (~(A25iu6 & Ppfpw6[10]));
assign Uqciu6 = (~(R05iu6 & D7fpw6[10]));
assign Jzuhu6 = (~(Irciu6 & Prciu6));
assign Prciu6 = (Wrciu6 & Dsciu6);
assign Dsciu6 = (~(HRDATA[9] & Pp7iu6));
assign Wrciu6 = (Ksciu6 & Rsciu6);
assign Rsciu6 = (~(Hrfpw6[9] & Uy4iu6));
assign Ksciu6 = (~(HRDATA[25] & Kq7iu6));
assign Irciu6 = (Ysciu6 & Ftciu6);
assign Ftciu6 = (~(A25iu6 & Ppfpw6[9]));
assign Ysciu6 = (~(R05iu6 & D7fpw6[9]));
assign Czuhu6 = (!Mtciu6);
assign Mtciu6 = (HREADY ? Auciu6 : Ttciu6);
assign Auciu6 = (~(Huciu6 & Ouciu6));
assign Ouciu6 = (Vuciu6 & Cvciu6);
assign Huciu6 = (HALTED & A2nhu6);
assign Vyuhu6 = (~(Jvciu6 & Qvciu6));
assign Qvciu6 = (~(Xvciu6 & Hv4iu6));
assign Hv4iu6 = (!Daohu6);
assign Xvciu6 = (~(HALTED & HREADY));
assign Jvciu6 = (Eh6iu6 | DBGRESTART);
assign Oyuhu6 = (~(Jw4iu6 & Ewciu6));
assign Ewciu6 = (~(Dhgpw6[4] & Lwciu6));
assign Lwciu6 = (~(Scbiu6 & H34iu6));
assign Jw4iu6 = (~(Swciu6 & EDBGRQ));
assign Swciu6 = (~(Zwciu6 | HALTED));
assign Hyuhu6 = (Wi7iu6 ? HWRITE : Gxciu6);
assign Wi7iu6 = (~(Bq6iu6 & Nxciu6));
assign Nxciu6 = (~(Uxciu6 & Byciu6));
assign Byciu6 = (~(Iyciu6 | Pyciu6));
assign Iyciu6 = (Wyciu6 | V0epw6);
assign Wyciu6 = (!Z18iu6);
assign Uxciu6 = (S18iu6 & Hy8iu6);
assign Bq6iu6 = (Dzciu6 | Kzciu6);
assign Dzciu6 = (~(Xg6iu6 & HREADY));
assign Gxciu6 = (Rzciu6 & Yzciu6);
assign Ayuhu6 = (~(F0diu6 & M0diu6));
assign M0diu6 = (~(Vbgpw6[30] & T0diu6));
assign T0diu6 = (~(HWDATA[30] & O59iu6));
assign F0diu6 = (~(V59iu6 & HWDATA[30]));
assign Txuhu6 = (Dv9iu6 ? R4gpw6[6] : HWDATA[30]);
assign Mxuhu6 = (~(A1diu6 & H1diu6));
assign H1diu6 = (~(Vbgpw6[29] & O1diu6));
assign O1diu6 = (~(HWDATA[29] & O59iu6));
assign A1diu6 = (~(V59iu6 & HWDATA[29]));
assign Fxuhu6 = (~(V1diu6 & C2diu6));
assign C2diu6 = (~(Vbgpw6[28] & J2diu6));
assign J2diu6 = (~(HWDATA[28] & O59iu6));
assign V1diu6 = (~(V59iu6 & HWDATA[28]));
assign Ywuhu6 = (~(Q2diu6 & X2diu6));
assign X2diu6 = (~(Vbgpw6[27] & E3diu6));
assign E3diu6 = (~(HWDATA[27] & O59iu6));
assign Q2diu6 = (~(V59iu6 & HWDATA[27]));
assign Rwuhu6 = (~(L3diu6 & S3diu6));
assign S3diu6 = (~(Vbgpw6[26] & Z3diu6));
assign Z3diu6 = (~(HWDATA[26] & O59iu6));
assign L3diu6 = (~(V59iu6 & HWDATA[26]));
assign Kwuhu6 = (~(G4diu6 & N4diu6));
assign N4diu6 = (~(Vbgpw6[25] & U4diu6));
assign U4diu6 = (~(HWDATA[25] & O59iu6));
assign G4diu6 = (~(V59iu6 & HWDATA[25]));
assign Dwuhu6 = (~(B5diu6 & I5diu6));
assign I5diu6 = (~(Vbgpw6[24] & P5diu6));
assign P5diu6 = (~(HWDATA[24] & O59iu6));
assign B5diu6 = (~(V59iu6 & HWDATA[24]));
assign Wvuhu6 = (~(W5diu6 & D6diu6));
assign D6diu6 = (~(Vbgpw6[23] & K6diu6));
assign K6diu6 = (~(HWDATA[23] & O59iu6));
assign W5diu6 = (~(V59iu6 & HWDATA[23]));
assign Pvuhu6 = (R6diu6 & Y6diu6);
assign Y6diu6 = (F7diu6 & M7diu6);
assign F7diu6 = (~(Drdpw6 & T7diu6));
assign R6diu6 = (IRQ[23] & A8diu6);
assign A8diu6 = (~(Tk7iu6 & H8diu6));
assign H8diu6 = (O8diu6 | Qg6iu6);
assign Ivuhu6 = (Dv9iu6 ? R4gpw6[5] : HWDATA[23]);
assign Bvuhu6 = (~(V8diu6 & C9diu6));
assign C9diu6 = (~(Vbgpw6[22] & J9diu6));
assign J9diu6 = (~(HWDATA[22] & O59iu6));
assign V8diu6 = (~(V59iu6 & HWDATA[22]));
assign Uuuhu6 = (Q9diu6 & X9diu6);
assign X9diu6 = (Eadiu6 & Ladiu6);
assign Eadiu6 = (~(Xndpw6 & Sadiu6));
assign Q9diu6 = (IRQ[22] & Zadiu6);
assign Zadiu6 = (~(Tk7iu6 & Gbdiu6));
assign Gbdiu6 = (Qg6iu6 | Nbdiu6);
assign Nuuhu6 = (Dv9iu6 ? R4gpw6[4] : HWDATA[22]);
assign Guuhu6 = (~(Ubdiu6 & Bcdiu6));
assign Bcdiu6 = (~(Vbgpw6[21] & Icdiu6));
assign Icdiu6 = (~(HWDATA[21] & O59iu6));
assign Ubdiu6 = (~(V59iu6 & HWDATA[21]));
assign Ztuhu6 = (Pcdiu6 & Wcdiu6);
assign Wcdiu6 = (Dddiu6 & Kddiu6);
assign Dddiu6 = (~(Rrdpw6 & Rddiu6));
assign Pcdiu6 = (IRQ[21] & Yddiu6);
assign Yddiu6 = (~(Tk7iu6 & Fediu6));
assign Fediu6 = (Mediu6 | Qg6iu6);
assign Stuhu6 = (~(Tediu6 & Afdiu6));
assign Afdiu6 = (~(Vbgpw6[20] & Hfdiu6));
assign Hfdiu6 = (~(HWDATA[20] & O59iu6));
assign Tediu6 = (~(V59iu6 & HWDATA[20]));
assign Ltuhu6 = (Ofdiu6 & Vfdiu6);
assign Vfdiu6 = (Cgdiu6 & Jgdiu6);
assign Cgdiu6 = (~(Yrdpw6 & Qgdiu6));
assign Ofdiu6 = (IRQ[20] & Xgdiu6);
assign Xgdiu6 = (~(Tk7iu6 & Ehdiu6));
assign Ehdiu6 = (Qg6iu6 | Lhdiu6);
assign Etuhu6 = (~(Shdiu6 & Zhdiu6));
assign Zhdiu6 = (~(Vbgpw6[19] & Gidiu6));
assign Gidiu6 = (~(HWDATA[19] & O59iu6));
assign Shdiu6 = (~(V59iu6 & HWDATA[19]));
assign Xsuhu6 = (Nidiu6 & Uidiu6);
assign Uidiu6 = (Bjdiu6 & Ijdiu6);
assign Bjdiu6 = (~(Msdpw6 & Pjdiu6));
assign Nidiu6 = (IRQ[19] & Wjdiu6);
assign Wjdiu6 = (~(Tk7iu6 & Dkdiu6));
assign Dkdiu6 = (Qg6iu6 | Kkdiu6);
assign Qsuhu6 = (~(Rkdiu6 & Ykdiu6));
assign Ykdiu6 = (~(Vbgpw6[18] & Fldiu6));
assign Fldiu6 = (~(HWDATA[18] & O59iu6));
assign Rkdiu6 = (~(V59iu6 & HWDATA[18]));
assign Jsuhu6 = (Mldiu6 & Tldiu6);
assign Tldiu6 = (Amdiu6 & Hmdiu6);
assign Amdiu6 = (~(Tsdpw6 & Omdiu6));
assign Mldiu6 = (IRQ[18] & Vmdiu6);
assign Vmdiu6 = (~(Tk7iu6 & Cndiu6));
assign Cndiu6 = (Qg6iu6 | Jndiu6);
assign Csuhu6 = (~(Qndiu6 & Xndiu6));
assign Xndiu6 = (~(Vbgpw6[17] & Eodiu6));
assign Eodiu6 = (~(HWDATA[17] & O59iu6));
assign Qndiu6 = (~(V59iu6 & HWDATA[17]));
assign Vruhu6 = (Lodiu6 & Sodiu6);
assign Sodiu6 = (Zodiu6 & Gpdiu6);
assign Zodiu6 = (~(Htdpw6 & Npdiu6));
assign Lodiu6 = (IRQ[17] & Updiu6);
assign Updiu6 = (~(Tk7iu6 & Bqdiu6));
assign Bqdiu6 = (Qg6iu6 | Iqdiu6);
assign Oruhu6 = (~(Pqdiu6 & Wqdiu6));
assign Wqdiu6 = (~(Vbgpw6[16] & Drdiu6));
assign Drdiu6 = (~(HWDATA[16] & O59iu6));
assign Pqdiu6 = (~(V59iu6 & HWDATA[16]));
assign Hruhu6 = (~(Krdiu6 & Rrdiu6));
assign Rrdiu6 = (~(Vbgpw6[15] & Yrdiu6));
assign Yrdiu6 = (~(Fsdiu6 & O59iu6));
assign Krdiu6 = (~(V59iu6 & Fsdiu6));
assign Aruhu6 = (Dv9iu6 ? R4gpw6[3] : Fsdiu6);
assign Tquhu6 = (~(Msdiu6 & Tsdiu6));
assign Tsdiu6 = (~(Vbgpw6[14] & Atdiu6));
assign Atdiu6 = (~(HWDATA[14] & O59iu6));
assign Msdiu6 = (~(V59iu6 & HWDATA[14]));
assign Mquhu6 = (Dv9iu6 ? R4gpw6[2] : HWDATA[14]);
assign Fquhu6 = (~(Htdiu6 & Otdiu6));
assign Otdiu6 = (~(Vbgpw6[13] & Vtdiu6));
assign Vtdiu6 = (~(HWDATA[13] & O59iu6));
assign Htdiu6 = (~(V59iu6 & HWDATA[13]));
assign Ypuhu6 = (~(Cudiu6 & Judiu6));
assign Judiu6 = (~(Vbgpw6[12] & Qudiu6));
assign Qudiu6 = (~(HWDATA[12] & O59iu6));
assign Cudiu6 = (~(V59iu6 & HWDATA[12]));
assign Rpuhu6 = (~(Xudiu6 & Evdiu6));
assign Evdiu6 = (~(Vbgpw6[11] & Lvdiu6));
assign Lvdiu6 = (~(HWDATA[11] & O59iu6));
assign Xudiu6 = (~(V59iu6 & HWDATA[11]));
assign Kpuhu6 = (~(Svdiu6 & Zvdiu6));
assign Zvdiu6 = (~(Vbgpw6[10] & Gwdiu6));
assign Gwdiu6 = (~(HWDATA[10] & O59iu6));
assign Svdiu6 = (~(V59iu6 & HWDATA[10]));
assign Dpuhu6 = (~(Nwdiu6 & Uwdiu6));
assign Uwdiu6 = (~(Vbgpw6[9] & Bxdiu6));
assign Bxdiu6 = (~(HWDATA[9] & O59iu6));
assign Nwdiu6 = (~(V59iu6 & HWDATA[9]));
assign Wouhu6 = (~(Ixdiu6 & Pxdiu6));
assign Pxdiu6 = (~(Vbgpw6[8] & Wxdiu6));
assign Wxdiu6 = (~(HWDATA[8] & O59iu6));
assign Ixdiu6 = (~(V59iu6 & HWDATA[8]));
assign Pouhu6 = (~(Dydiu6 & Kydiu6));
assign Kydiu6 = (~(Vbgpw6[7] & Rydiu6));
assign Rydiu6 = (~(HWDATA[7] & O59iu6));
assign Dydiu6 = (~(V59iu6 & HWDATA[7]));
assign Iouhu6 = (Dv9iu6 ? R4gpw6[1] : HWDATA[7]);
assign Bouhu6 = (~(Yydiu6 & Fzdiu6));
assign Fzdiu6 = (~(Vbgpw6[6] & Mzdiu6));
assign Mzdiu6 = (~(HWDATA[6] & O59iu6));
assign Yydiu6 = (~(V59iu6 & HWDATA[6]));
assign Unuhu6 = (Dv9iu6 ? R4gpw6[0] : HWDATA[6]);
assign Dv9iu6 = (~(Tzdiu6 & Npdhu6));
assign Nnuhu6 = (~(A0eiu6 & H0eiu6));
assign H0eiu6 = (~(Vbgpw6[5] & O0eiu6));
assign O0eiu6 = (~(HWDATA[5] & O59iu6));
assign A0eiu6 = (~(V59iu6 & HWDATA[5]));
assign Gnuhu6 = (~(V0eiu6 & C1eiu6));
assign C1eiu6 = (~(Vbgpw6[4] & J1eiu6));
assign J1eiu6 = (~(HWDATA[4] & O59iu6));
assign V0eiu6 = (~(V59iu6 & HWDATA[4]));
assign Zmuhu6 = (~(Q1eiu6 & X1eiu6));
assign X1eiu6 = (~(Vbgpw6[3] & E2eiu6));
assign E2eiu6 = (~(HWDATA[3] & O59iu6));
assign Q1eiu6 = (~(V59iu6 & HWDATA[3]));
assign Smuhu6 = (~(L2eiu6 & S2eiu6));
assign S2eiu6 = (~(Vbgpw6[2] & Z2eiu6));
assign Z2eiu6 = (~(G3eiu6 & O59iu6));
assign L2eiu6 = (~(V59iu6 & G3eiu6));
assign Lmuhu6 = (~(N3eiu6 & U3eiu6));
assign U3eiu6 = (~(Vbgpw6[1] & B4eiu6));
assign B4eiu6 = (~(I4eiu6 & O59iu6));
assign O59iu6 = (V59iu6 | P4eiu6);
assign P4eiu6 = (W4eiu6 & D5eiu6);
assign W4eiu6 = (Npdhu6 & K5eiu6);
assign N3eiu6 = (~(V59iu6 & I4eiu6));
assign V59iu6 = (Yzciu6 & K5eiu6);
assign Emuhu6 = (R5eiu6 ? Bxghu6 : HWDATA[0]);
assign Xluhu6 = (R5eiu6 ? Ftghu6 : G3eiu6);
assign Qluhu6 = (R5eiu6 ? Dvghu6 : I4eiu6);
assign R5eiu6 = (~(Y5eiu6 & Npdhu6));
assign Jluhu6 = (F6eiu6 ? Bagpw6[0] : HWDATA[0]);
assign Cluhu6 = (F6eiu6 ? Bagpw6[23] : HWDATA[23]);
assign Vkuhu6 = (F6eiu6 ? Bagpw6[22] : HWDATA[22]);
assign Okuhu6 = (F6eiu6 ? Bagpw6[21] : HWDATA[21]);
assign Hkuhu6 = (F6eiu6 ? Bagpw6[20] : HWDATA[20]);
assign Akuhu6 = (F6eiu6 ? Bagpw6[19] : HWDATA[19]);
assign Tjuhu6 = (F6eiu6 ? Bagpw6[18] : HWDATA[18]);
assign Mjuhu6 = (F6eiu6 ? Bagpw6[17] : HWDATA[17]);
assign Fjuhu6 = (F6eiu6 ? Bagpw6[16] : HWDATA[16]);
assign Yiuhu6 = (F6eiu6 ? Bagpw6[15] : Fsdiu6);
assign Riuhu6 = (F6eiu6 ? Bagpw6[14] : HWDATA[14]);
assign Kiuhu6 = (F6eiu6 ? Bagpw6[13] : HWDATA[13]);
assign Diuhu6 = (F6eiu6 ? Bagpw6[12] : HWDATA[12]);
assign Whuhu6 = (F6eiu6 ? Bagpw6[11] : HWDATA[11]);
assign Phuhu6 = (F6eiu6 ? Bagpw6[10] : HWDATA[10]);
assign Ihuhu6 = (F6eiu6 ? Bagpw6[9] : HWDATA[9]);
assign Bhuhu6 = (F6eiu6 ? Bagpw6[8] : HWDATA[8]);
assign Uguhu6 = (F6eiu6 ? Bagpw6[7] : HWDATA[7]);
assign Nguhu6 = (F6eiu6 ? Bagpw6[6] : HWDATA[6]);
assign Gguhu6 = (F6eiu6 ? Bagpw6[5] : HWDATA[5]);
assign Zfuhu6 = (F6eiu6 ? Bagpw6[4] : HWDATA[4]);
assign Sfuhu6 = (F6eiu6 ? Bagpw6[3] : HWDATA[3]);
assign Lfuhu6 = (F6eiu6 ? Bagpw6[2] : G3eiu6);
assign Efuhu6 = (F6eiu6 ? Bagpw6[1] : I4eiu6);
assign F6eiu6 = (~(M6eiu6 & Npdhu6));
assign Xeuhu6 = (~(T6eiu6 & A7eiu6));
assign A7eiu6 = (H7eiu6 | O7eiu6);
assign T6eiu6 = (V7eiu6 & C8eiu6);
assign C8eiu6 = (~(L6gpw6[0] & J8eiu6));
assign V7eiu6 = (~(Q8eiu6 & Bagpw6[0]));
assign Qeuhu6 = (~(X8eiu6 & E9eiu6));
assign E9eiu6 = (~(L9eiu6 & Tzfpw6[1]));
assign X8eiu6 = (S9eiu6 & Z9eiu6);
assign Z9eiu6 = (~(L6gpw6[1] & J8eiu6));
assign S9eiu6 = (~(Q8eiu6 & Bagpw6[1]));
assign Jeuhu6 = (~(Gaeiu6 & Naeiu6));
assign Naeiu6 = (~(L9eiu6 & Tzfpw6[2]));
assign Gaeiu6 = (Uaeiu6 & Bbeiu6);
assign Bbeiu6 = (~(L6gpw6[2] & J8eiu6));
assign Uaeiu6 = (~(Q8eiu6 & Bagpw6[2]));
assign Ceuhu6 = (~(Ibeiu6 & Pbeiu6));
assign Pbeiu6 = (~(Tzfpw6[3] & L9eiu6));
assign Ibeiu6 = (Wbeiu6 & Dceiu6);
assign Dceiu6 = (~(L6gpw6[3] & J8eiu6));
assign Wbeiu6 = (~(Q8eiu6 & Bagpw6[3]));
assign Vduhu6 = (~(Kceiu6 & Rceiu6));
assign Rceiu6 = (~(L9eiu6 & Tzfpw6[4]));
assign Kceiu6 = (Yceiu6 & Fdeiu6);
assign Fdeiu6 = (~(L6gpw6[4] & J8eiu6));
assign Yceiu6 = (~(Q8eiu6 & Bagpw6[4]));
assign Oduhu6 = (~(Mdeiu6 & Tdeiu6));
assign Tdeiu6 = (~(L9eiu6 & Tzfpw6[5]));
assign Mdeiu6 = (Aeeiu6 & Heeiu6);
assign Heeiu6 = (~(L6gpw6[5] & J8eiu6));
assign Aeeiu6 = (~(Q8eiu6 & Bagpw6[5]));
assign Hduhu6 = (~(Oeeiu6 & Veeiu6));
assign Veeiu6 = (~(L9eiu6 & Tzfpw6[6]));
assign Oeeiu6 = (Cfeiu6 & Jfeiu6);
assign Jfeiu6 = (~(L6gpw6[6] & J8eiu6));
assign Cfeiu6 = (~(Q8eiu6 & Bagpw6[6]));
assign Aduhu6 = (~(Qfeiu6 & Xfeiu6));
assign Xfeiu6 = (~(L9eiu6 & Tzfpw6[7]));
assign Qfeiu6 = (Egeiu6 & Lgeiu6);
assign Lgeiu6 = (~(L6gpw6[7] & J8eiu6));
assign Egeiu6 = (~(Q8eiu6 & Bagpw6[7]));
assign Tcuhu6 = (~(Sgeiu6 & Zgeiu6));
assign Zgeiu6 = (~(L9eiu6 & Tzfpw6[8]));
assign Sgeiu6 = (Gheiu6 & Nheiu6);
assign Nheiu6 = (~(L6gpw6[8] & J8eiu6));
assign Gheiu6 = (~(Q8eiu6 & Bagpw6[8]));
assign Mcuhu6 = (~(Uheiu6 & Bieiu6));
assign Bieiu6 = (~(L9eiu6 & Tzfpw6[9]));
assign Uheiu6 = (Iieiu6 & Pieiu6);
assign Pieiu6 = (~(L6gpw6[9] & J8eiu6));
assign Iieiu6 = (~(Q8eiu6 & Bagpw6[9]));
assign Fcuhu6 = (~(Wieiu6 & Djeiu6));
assign Djeiu6 = (~(L9eiu6 & Tzfpw6[10]));
assign Wieiu6 = (Kjeiu6 & Rjeiu6);
assign Rjeiu6 = (~(L6gpw6[10] & J8eiu6));
assign Kjeiu6 = (~(Q8eiu6 & Bagpw6[10]));
assign Ybuhu6 = (~(Yjeiu6 & Fkeiu6));
assign Fkeiu6 = (~(Tzfpw6[11] & L9eiu6));
assign Yjeiu6 = (Mkeiu6 & Tkeiu6);
assign Tkeiu6 = (~(L6gpw6[11] & J8eiu6));
assign Mkeiu6 = (~(Q8eiu6 & Bagpw6[11]));
assign Rbuhu6 = (~(Aleiu6 & Hleiu6));
assign Hleiu6 = (~(L9eiu6 & Tzfpw6[12]));
assign Aleiu6 = (Oleiu6 & Vleiu6);
assign Vleiu6 = (~(L6gpw6[12] & J8eiu6));
assign Oleiu6 = (~(Q8eiu6 & Bagpw6[12]));
assign Kbuhu6 = (~(Cmeiu6 & Jmeiu6));
assign Jmeiu6 = (~(L9eiu6 & Tzfpw6[13]));
assign Cmeiu6 = (Qmeiu6 & Xmeiu6);
assign Xmeiu6 = (~(L6gpw6[13] & J8eiu6));
assign Qmeiu6 = (~(Q8eiu6 & Bagpw6[13]));
assign Dbuhu6 = (~(Eneiu6 & Lneiu6));
assign Lneiu6 = (~(L9eiu6 & Tzfpw6[14]));
assign Eneiu6 = (Sneiu6 & Zneiu6);
assign Zneiu6 = (~(L6gpw6[14] & J8eiu6));
assign Sneiu6 = (~(Q8eiu6 & Bagpw6[14]));
assign Wauhu6 = (~(Goeiu6 & Noeiu6));
assign Noeiu6 = (~(L9eiu6 & Tzfpw6[15]));
assign Goeiu6 = (Uoeiu6 & Bpeiu6);
assign Bpeiu6 = (~(L6gpw6[15] & J8eiu6));
assign Uoeiu6 = (~(Q8eiu6 & Bagpw6[15]));
assign Pauhu6 = (~(Ipeiu6 & Ppeiu6));
assign Ppeiu6 = (~(L9eiu6 & Tzfpw6[16]));
assign Ipeiu6 = (Wpeiu6 & Dqeiu6);
assign Dqeiu6 = (~(L6gpw6[16] & J8eiu6));
assign Wpeiu6 = (~(Q8eiu6 & Bagpw6[16]));
assign Iauhu6 = (~(Kqeiu6 & Rqeiu6));
assign Rqeiu6 = (~(L9eiu6 & Tzfpw6[17]));
assign Kqeiu6 = (Yqeiu6 & Freiu6);
assign Freiu6 = (~(L6gpw6[17] & J8eiu6));
assign Yqeiu6 = (~(Q8eiu6 & Bagpw6[17]));
assign Bauhu6 = (~(Mreiu6 & Treiu6));
assign Treiu6 = (~(L9eiu6 & Tzfpw6[18]));
assign Mreiu6 = (Aseiu6 & Hseiu6);
assign Hseiu6 = (~(L6gpw6[18] & J8eiu6));
assign Aseiu6 = (~(Q8eiu6 & Bagpw6[18]));
assign U9uhu6 = (~(Oseiu6 & Vseiu6));
assign Vseiu6 = (~(Tzfpw6[19] & L9eiu6));
assign Oseiu6 = (Cteiu6 & Jteiu6);
assign Jteiu6 = (~(L6gpw6[19] & J8eiu6));
assign Cteiu6 = (~(Q8eiu6 & Bagpw6[19]));
assign N9uhu6 = (~(Qteiu6 & Xteiu6));
assign Xteiu6 = (~(L9eiu6 & Tzfpw6[20]));
assign Qteiu6 = (Eueiu6 & Lueiu6);
assign Lueiu6 = (~(L6gpw6[20] & J8eiu6));
assign Eueiu6 = (~(Q8eiu6 & Bagpw6[20]));
assign G9uhu6 = (~(Sueiu6 & Zueiu6));
assign Zueiu6 = (~(L9eiu6 & Tzfpw6[21]));
assign Sueiu6 = (Gveiu6 & Nveiu6);
assign Nveiu6 = (~(L6gpw6[21] & J8eiu6));
assign Gveiu6 = (~(Q8eiu6 & Bagpw6[21]));
assign Z8uhu6 = (~(Uveiu6 & Bweiu6));
assign Bweiu6 = (~(L9eiu6 & Tzfpw6[22]));
assign Uveiu6 = (Iweiu6 & Pweiu6);
assign Pweiu6 = (~(L6gpw6[22] & J8eiu6));
assign Iweiu6 = (~(Q8eiu6 & Bagpw6[22]));
assign S8uhu6 = (~(Wweiu6 & Dxeiu6));
assign Dxeiu6 = (~(L9eiu6 & Tzfpw6[23]));
assign Wweiu6 = (Kxeiu6 & Rxeiu6);
assign Rxeiu6 = (~(L6gpw6[23] & J8eiu6));
assign J8eiu6 = (Yxeiu6 & Fyeiu6);
assign Yxeiu6 = (~(L9eiu6 | Myeiu6));
assign Kxeiu6 = (~(Q8eiu6 & Bagpw6[23]));
assign Q8eiu6 = (~(Tyeiu6 | Fyeiu6));
assign Fyeiu6 = (~(Azeiu6 & O7eiu6));
assign O7eiu6 = (!Tzfpw6[0]);
assign Tyeiu6 = (~(H7eiu6 & Hzeiu6));
assign H7eiu6 = (!L9eiu6);
assign L9eiu6 = (~(Ozeiu6 | Myeiu6));
assign Myeiu6 = (!Hzeiu6);
assign L8uhu6 = (Vzeiu6 ? R4gpw6[56] : HWDATA[6]);
assign E8uhu6 = (Vzeiu6 ? R4gpw6[57] : HWDATA[7]);
assign X7uhu6 = (Vzeiu6 ? R4gpw6[58] : HWDATA[14]);
assign Q7uhu6 = (Vzeiu6 ? R4gpw6[59] : Fsdiu6);
assign J7uhu6 = (Vzeiu6 ? R4gpw6[60] : HWDATA[22]);
assign C7uhu6 = (Vzeiu6 ? R4gpw6[61] : HWDATA[23]);
assign V6uhu6 = (Vzeiu6 ? R4gpw6[62] : HWDATA[30]);
assign O6uhu6 = (Vzeiu6 ? R4gpw6[63] : HWDATA[31]);
assign Vzeiu6 = (~(C0fiu6 & Npdhu6));
assign H6uhu6 = (J0fiu6 ? R4gpw6[48] : HWDATA[6]);
assign A6uhu6 = (J0fiu6 ? R4gpw6[49] : HWDATA[7]);
assign T5uhu6 = (J0fiu6 ? R4gpw6[50] : HWDATA[14]);
assign M5uhu6 = (J0fiu6 ? R4gpw6[51] : Fsdiu6);
assign F5uhu6 = (J0fiu6 ? R4gpw6[52] : HWDATA[22]);
assign Y4uhu6 = (J0fiu6 ? R4gpw6[53] : HWDATA[23]);
assign R4uhu6 = (J0fiu6 ? R4gpw6[54] : HWDATA[30]);
assign K4uhu6 = (J0fiu6 ? R4gpw6[55] : HWDATA[31]);
assign J0fiu6 = (~(Q0fiu6 & Npdhu6));
assign D4uhu6 = (X0fiu6 ? R4gpw6[40] : HWDATA[6]);
assign W3uhu6 = (X0fiu6 ? R4gpw6[41] : HWDATA[7]);
assign P3uhu6 = (X0fiu6 ? R4gpw6[42] : HWDATA[14]);
assign I3uhu6 = (X0fiu6 ? R4gpw6[43] : Fsdiu6);
assign B3uhu6 = (X0fiu6 ? R4gpw6[44] : HWDATA[22]);
assign U2uhu6 = (X0fiu6 ? R4gpw6[45] : HWDATA[23]);
assign N2uhu6 = (X0fiu6 ? R4gpw6[46] : HWDATA[30]);
assign G2uhu6 = (X0fiu6 ? R4gpw6[47] : HWDATA[31]);
assign X0fiu6 = (~(E1fiu6 & Npdhu6));
assign Z1uhu6 = (L1fiu6 ? R4gpw6[32] : HWDATA[6]);
assign S1uhu6 = (L1fiu6 ? R4gpw6[33] : HWDATA[7]);
assign L1uhu6 = (L1fiu6 ? R4gpw6[34] : HWDATA[14]);
assign E1uhu6 = (L1fiu6 ? R4gpw6[35] : Fsdiu6);
assign X0uhu6 = (L1fiu6 ? R4gpw6[36] : HWDATA[22]);
assign Q0uhu6 = (L1fiu6 ? R4gpw6[37] : HWDATA[23]);
assign J0uhu6 = (L1fiu6 ? R4gpw6[38] : HWDATA[30]);
assign C0uhu6 = (L1fiu6 ? R4gpw6[39] : HWDATA[31]);
assign L1fiu6 = (~(S1fiu6 & Npdhu6));
assign Vzthu6 = (Z1fiu6 ? R4gpw6[24] : HWDATA[6]);
assign Ozthu6 = (Z1fiu6 ? R4gpw6[25] : HWDATA[7]);
assign Hzthu6 = (Z1fiu6 ? R4gpw6[26] : HWDATA[14]);
assign Azthu6 = (Z1fiu6 ? R4gpw6[27] : Fsdiu6);
assign Tythu6 = (Z1fiu6 ? R4gpw6[28] : HWDATA[22]);
assign Mythu6 = (Z1fiu6 ? R4gpw6[29] : HWDATA[23]);
assign Fythu6 = (Z1fiu6 ? R4gpw6[30] : HWDATA[30]);
assign Yxthu6 = (Z1fiu6 ? R4gpw6[31] : HWDATA[31]);
assign Z1fiu6 = (~(G2fiu6 & Npdhu6));
assign Rxthu6 = (N2fiu6 ? R4gpw6[16] : HWDATA[6]);
assign Kxthu6 = (N2fiu6 ? R4gpw6[17] : HWDATA[7]);
assign Dxthu6 = (N2fiu6 ? R4gpw6[18] : HWDATA[14]);
assign Wwthu6 = (N2fiu6 ? R4gpw6[19] : Fsdiu6);
assign Pwthu6 = (N2fiu6 ? R4gpw6[20] : HWDATA[22]);
assign Iwthu6 = (N2fiu6 ? R4gpw6[21] : HWDATA[23]);
assign Bwthu6 = (N2fiu6 ? R4gpw6[22] : HWDATA[30]);
assign Uvthu6 = (N2fiu6 ? R4gpw6[23] : HWDATA[31]);
assign N2fiu6 = (~(U2fiu6 & Npdhu6));
assign Nvthu6 = (B3fiu6 ? R4gpw6[8] : HWDATA[6]);
assign Gvthu6 = (B3fiu6 ? R4gpw6[9] : HWDATA[7]);
assign Zuthu6 = (B3fiu6 ? R4gpw6[10] : HWDATA[14]);
assign Suthu6 = (B3fiu6 ? R4gpw6[11] : Fsdiu6);
assign Luthu6 = (B3fiu6 ? R4gpw6[12] : HWDATA[22]);
assign Euthu6 = (B3fiu6 ? R4gpw6[13] : HWDATA[23]);
assign Xtthu6 = (B3fiu6 ? R4gpw6[14] : HWDATA[30]);
assign Qtthu6 = (B3fiu6 ? R4gpw6[15] : HWDATA[31]);
assign B3fiu6 = (~(I3fiu6 & Npdhu6));
assign Jtthu6 = (P3fiu6 ? Gfghu6 : HWDATA[4]);
assign Ctthu6 = (~(W3fiu6 & D4fiu6));
assign D4fiu6 = (~(vis_ipsr_o[4] & F8ciu6));
assign W3fiu6 = (K4fiu6 & R4fiu6);
assign R4fiu6 = (~(Xibiu6 & Ppfpw6[4]));
assign K4fiu6 = (Ejbiu6 | Y4fiu6);
assign Vsthu6 = (F5fiu6 & M5fiu6);
assign M5fiu6 = (T5fiu6 & A6fiu6);
assign T5fiu6 = (~(Zodpw6 & H6fiu6));
assign F5fiu6 = (IRQ[7] & O6fiu6);
assign O6fiu6 = (~(Tk7iu6 & V6fiu6));
assign V6fiu6 = (Qg6iu6 | C7fiu6);
assign Osthu6 = (J7fiu6 & Q7fiu6);
assign Q7fiu6 = (X7fiu6 & E8fiu6);
assign X7fiu6 = (~(Lodpw6 & L8fiu6));
assign J7fiu6 = (IRQ[6] & S8fiu6);
assign S8fiu6 = (~(Tk7iu6 & Z8fiu6));
assign Z8fiu6 = (G9fiu6 | Qg6iu6);
assign Hsthu6 = (N9fiu6 & U9fiu6);
assign U9fiu6 = (Bafiu6 & Iafiu6);
assign Bafiu6 = (~(Gpdpw6 & Pafiu6));
assign N9fiu6 = (IRQ[5] & Wafiu6);
assign Wafiu6 = (~(Tk7iu6 & Dbfiu6));
assign Dbfiu6 = (Kbfiu6 | Qg6iu6);
assign Asthu6 = (Rbfiu6 & Ybfiu6);
assign Ybfiu6 = (Fcfiu6 & Mcfiu6);
assign Fcfiu6 = (~(Qndpw6 & Tcfiu6));
assign Rbfiu6 = (IRQ[4] & Adfiu6);
assign Adfiu6 = (~(Tk7iu6 & Hdfiu6));
assign Hdfiu6 = (Qg6iu6 | Odfiu6);
assign Trthu6 = (Vdfiu6 & Cefiu6);
assign Cefiu6 = (Jefiu6 & Qefiu6);
assign Jefiu6 = (~(Jndpw6 & Xefiu6));
assign Vdfiu6 = (IRQ[3] & Effiu6);
assign Effiu6 = (~(Tk7iu6 & Lffiu6));
assign Lffiu6 = (Sffiu6 | Qg6iu6);
assign Mrthu6 = (~(Zffiu6 & Ggfiu6));
assign Ggfiu6 = (Ngfiu6 | Cibiu6);
assign Zffiu6 = (Ugfiu6 & Bhfiu6);
assign Bhfiu6 = (~(Xibiu6 & Ppfpw6[3]));
assign Xibiu6 = (Ihfiu6 & Phfiu6);
assign Phfiu6 = (~(Qaciu6 | Qg6iu6));
assign Qaciu6 = (~(Whfiu6 | Difiu6));
assign Ihfiu6 = (Cibiu6 & Ivfhu6);
assign Ugfiu6 = (Ejbiu6 | Kifiu6);
assign Ejbiu6 = (~(Rifiu6 & Cibiu6));
assign Cibiu6 = (!F8ciu6);
assign F8ciu6 = (~(HREADY & Yifiu6));
assign Yifiu6 = (~(Uzaiu6 & Fjfiu6));
assign Rifiu6 = (~(Mjfiu6 | Qg6iu6));
assign Frthu6 = (~(Xw4iu6 & Tjfiu6));
assign Tjfiu6 = (~(Dhgpw6[3] & Akfiu6));
assign Akfiu6 = (~(Scbiu6 & Df4iu6));
assign Xw4iu6 = (~(Jehhu6 & Hkfiu6));
assign Hkfiu6 = (~(Okfiu6 & Vkfiu6));
assign Vkfiu6 = (~(S3hhu6 & Ptaiu6));
assign Ptaiu6 = (M2biu6 & Clfiu6);
assign Okfiu6 = (~(H2hhu6 & Mu4iu6));
assign Yqthu6 = (Jlfiu6 & Qlfiu6);
assign Qlfiu6 = (Xlfiu6 & Jg6iu6);
assign Jg6iu6 = (~(Ch5iu6 & HWDATA[31]));
assign Xlfiu6 = (~(Evdpw6 & Af6iu6));
assign Af6iu6 = (Emfiu6 | Sb5iu6);
assign Jlfiu6 = (NMI & Lmfiu6);
assign Lmfiu6 = (~(Tk7iu6 & Smfiu6));
assign Smfiu6 = (Qg6iu6 | Zmfiu6);
assign Rqthu6 = (~(Gnfiu6 & Nnfiu6));
assign Nnfiu6 = (Unfiu6 | Bofiu6);
assign Bofiu6 = (L3ehu6 ? Ruaiu6 : Iofiu6);
assign Iofiu6 = (~(Uzaiu6 & Zmfiu6));
assign Unfiu6 = (~(F2biu6 & Sbghu6));
assign Gnfiu6 = (~(Jydhu6 & T2biu6));
assign T2biu6 = (~(HREADY & Pofiu6));
assign Pofiu6 = (Wofiu6 | C0ehu6);
assign Kqthu6 = (Dpfiu6 & Kpfiu6);
assign Kpfiu6 = (Rpfiu6 & Ypfiu6);
assign Rpfiu6 = (~(Bqdpw6 & Fqfiu6));
assign Dpfiu6 = (IRQ[28] & Mqfiu6);
assign Mqfiu6 = (~(Tk7iu6 & Tqfiu6));
assign Tqfiu6 = (Qg6iu6 | Arfiu6);
assign Dqthu6 = (Hrfiu6 & Orfiu6);
assign Orfiu6 = (Vrfiu6 & Csfiu6);
assign Vrfiu6 = (~(Iqdpw6 & Jsfiu6));
assign Hrfiu6 = (IRQ[27] & Qsfiu6);
assign Qsfiu6 = (~(Tk7iu6 & Xsfiu6));
assign Xsfiu6 = (Etfiu6 | Qg6iu6);
assign Wpthu6 = (Ltfiu6 & Stfiu6);
assign Stfiu6 = (Ztfiu6 & Gufiu6);
assign Ztfiu6 = (~(Pqdpw6 & Nufiu6));
assign Ltfiu6 = (IRQ[26] & Uufiu6);
assign Uufiu6 = (~(Tk7iu6 & Bvfiu6));
assign Bvfiu6 = (Ivfiu6 | Qg6iu6);
assign Ppthu6 = (Pvfiu6 & Wvfiu6);
assign Wvfiu6 = (Dwfiu6 & Fe6iu6);
assign Fe6iu6 = (~(Kwfiu6 & HWDATA[25]));
assign Dwfiu6 = (~(Krdpw6 & Wc6iu6));
assign Wc6iu6 = (Sb5iu6 | Rwfiu6);
assign Pvfiu6 = (IRQ[25] & Ywfiu6);
assign Ywfiu6 = (~(Tk7iu6 & Fxfiu6));
assign Fxfiu6 = (Mxfiu6 | Qg6iu6);
assign Ipthu6 = (Txfiu6 & Ayfiu6);
assign Ayfiu6 = (Hyfiu6 & Nb6iu6);
assign Nb6iu6 = (~(Kwfiu6 & HWDATA[24]));
assign Hyfiu6 = (~(Wqdpw6 & Ea6iu6));
assign Ea6iu6 = (Sb5iu6 | Oyfiu6);
assign Txfiu6 = (IRQ[24] & Vyfiu6);
assign Vyfiu6 = (~(Tk7iu6 & Czfiu6));
assign Czfiu6 = (Qg6iu6 | Jzfiu6);
assign Bpthu6 = (Qzfiu6 & Xzfiu6);
assign Xzfiu6 = (E0giu6 & L0giu6);
assign E0giu6 = (~(Lvdpw6 & S0giu6));
assign Qzfiu6 = (IRQ[15] & Z0giu6);
assign Z0giu6 = (~(Tk7iu6 & G1giu6));
assign G1giu6 = (N1giu6 | Qg6iu6);
assign Uothu6 = (U1giu6 & B2giu6);
assign B2giu6 = (I2giu6 & P2giu6);
assign I2giu6 = (~(Otdpw6 & W2giu6));
assign U1giu6 = (IRQ[14] & D3giu6);
assign D3giu6 = (~(Tk7iu6 & K3giu6));
assign K3giu6 = (R3giu6 | Qg6iu6);
assign Nothu6 = (Y3giu6 & F4giu6);
assign F4giu6 = (M4giu6 & T4giu6);
assign M4giu6 = (~(Vtdpw6 & A5giu6));
assign Y3giu6 = (IRQ[13] & H5giu6);
assign H5giu6 = (~(Tk7iu6 & O5giu6));
assign O5giu6 = (Qg6iu6 | V5giu6);
assign Gothu6 = (C6giu6 & J6giu6);
assign J6giu6 = (Q6giu6 & X6giu6);
assign Q6giu6 = (~(Qudpw6 & E7giu6));
assign C6giu6 = (IRQ[12] & L7giu6);
assign L7giu6 = (~(Tk7iu6 & S7giu6));
assign S7giu6 = (Qg6iu6 | Z7giu6);
assign Znthu6 = (G8giu6 & N8giu6);
assign N8giu6 = (U8giu6 & B9giu6);
assign U8giu6 = (~(Cudpw6 & I9giu6));
assign G8giu6 = (IRQ[11] & P9giu6);
assign P9giu6 = (~(Tk7iu6 & W9giu6));
assign W9giu6 = (Dagiu6 | Qg6iu6);
assign Snthu6 = (Kagiu6 & Ragiu6);
assign Ragiu6 = (Yagiu6 & Fbgiu6);
assign Yagiu6 = (~(Judpw6 & Mbgiu6));
assign Kagiu6 = (IRQ[10] & Tbgiu6);
assign Tbgiu6 = (~(Tk7iu6 & Acgiu6));
assign Acgiu6 = (Hcgiu6 | Qg6iu6);
assign Lnthu6 = (Ocgiu6 & Vcgiu6);
assign Vcgiu6 = (Cdgiu6 & J96iu6);
assign J96iu6 = (~(Kwfiu6 & HWDATA[9]));
assign Cdgiu6 = (~(Cndpw6 & A86iu6));
assign A86iu6 = (Sb5iu6 | Jdgiu6);
assign Ocgiu6 = (IRQ[9] & Qdgiu6);
assign Qdgiu6 = (~(Tk7iu6 & Xdgiu6));
assign Xdgiu6 = (Eegiu6 | Qg6iu6);
assign Enthu6 = (Legiu6 & Segiu6);
assign Segiu6 = (Zegiu6 & W56iu6);
assign W56iu6 = (~(Kwfiu6 & HWDATA[8]));
assign Zegiu6 = (~(Sodpw6 & N46iu6));
assign N46iu6 = (Sb5iu6 | Gfgiu6);
assign Legiu6 = (IRQ[8] & Nfgiu6);
assign Nfgiu6 = (~(Tk7iu6 & Ufgiu6));
assign Ufgiu6 = (Qg6iu6 | Bggiu6);
assign Xmthu6 = (~(Iggiu6 & Pggiu6));
assign Pggiu6 = (~(Ch5iu6 & HWDATA[28]));
assign Iggiu6 = (~(Wggiu6 & Ikghu6));
assign Wggiu6 = (Dhgiu6 & Khgiu6);
assign Khgiu6 = (~(Ch5iu6 & HWDATA[27]));
assign Dhgiu6 = (~(Clfiu6 & Rhgiu6));
assign Qmthu6 = (~(Ag5iu6 & Yhgiu6));
assign Yhgiu6 = (~(Figiu6 & Yyghu6));
assign Figiu6 = (Migiu6 & Tigiu6);
assign Tigiu6 = (~(Ch5iu6 & HWDATA[25]));
assign Migiu6 = (~(Clfiu6 & Ajgiu6));
assign Ag5iu6 = (Hjgiu6 & Ojgiu6);
assign Ojgiu6 = (~(Vjgiu6 & Ckgiu6));
assign Vjgiu6 = (Dvghu6 & Tzfpw6[0]);
assign Hjgiu6 = (~(Ch5iu6 & HWDATA[26]));
assign Ch5iu6 = (~(Jkgiu6 | Qkgiu6));
assign Jmthu6 = (Xkgiu6 & Elgiu6);
assign Elgiu6 = (Llgiu6 & Slgiu6);
assign Llgiu6 = (~(Eodpw6 & Zlgiu6));
assign Xkgiu6 = (IRQ[2] & Gmgiu6);
assign Gmgiu6 = (~(Tk7iu6 & Nmgiu6));
assign Nmgiu6 = (Qg6iu6 | Umgiu6);
assign Cmthu6 = (Bngiu6 & Ingiu6);
assign Ingiu6 = (Pngiu6 & Wngiu6);
assign Pngiu6 = (~(Fsdpw6 & Dogiu6));
assign Bngiu6 = (IRQ[1] & Kogiu6);
assign Kogiu6 = (~(Tk7iu6 & Rogiu6));
assign Rogiu6 = (Qg6iu6 | Yogiu6);
assign Vlthu6 = (P3fiu6 ? Qqdhu6 : I4eiu6);
assign Olthu6 = (P3fiu6 ? Ndghu6 : G3eiu6);
assign P3fiu6 = (~(Fpgiu6 & Npdhu6));
assign Hlthu6 = (Mpgiu6 ? B3gpw6[0] : HWDATA[30]);
assign Althu6 = (Mpgiu6 ? B3gpw6[1] : HWDATA[31]);
assign Mpgiu6 = (Tpgiu6 | Jkgiu6);
assign Tkthu6 = (Aqgiu6 ? L1gpw6[0] : HWDATA[22]);
assign Mkthu6 = (Aqgiu6 ? L1gpw6[1] : HWDATA[23]);
assign Fkthu6 = (Aqgiu6 ? H8gpw6[0] : HWDATA[30]);
assign Yjthu6 = (Aqgiu6 ? H8gpw6[1] : HWDATA[31]);
assign Aqgiu6 = (~(Hqgiu6 & Npdhu6));
assign Rjthu6 = (~(Qh5iu6 & Oqgiu6));
assign Oqgiu6 = (~(Vqgiu6 & Zlghu6));
assign Vqgiu6 = (Crgiu6 & Jrgiu6);
assign Jrgiu6 = (~(Clfiu6 & Qrgiu6));
assign Crgiu6 = (~(Xrgiu6 & Npdhu6));
assign Qh5iu6 = (Esgiu6 & Lsgiu6);
assign Lsgiu6 = (~(P0biu6 & Ssgiu6));
assign Ssgiu6 = (~(I0biu6 & Zsgiu6));
assign Zsgiu6 = (Gtgiu6 | Ntgiu6);
assign I0biu6 = (~(Utgiu6 & Bugiu6));
assign Bugiu6 = (~(Ae0iu6 | Cyfpw6[4]));
assign Utgiu6 = (Iugiu6 & Pugiu6);
assign Esgiu6 = (~(Xrgiu6 & Fsdiu6));
assign Kjthu6 = (~(Wugiu6 & Dvgiu6));
assign Dvgiu6 = (~(Kvgiu6 & Krghu6));
assign Kvgiu6 = (Rvgiu6 & Hzeiu6);
assign Hzeiu6 = (~(Yvgiu6 & Npdhu6));
assign Rvgiu6 = (~(Fwgiu6 & Y5eiu6));
assign Fwgiu6 = (Ur4iu6 & Jkgiu6);
assign Wugiu6 = (~(Ckgiu6 & Tzfpw6[0]));
assign Ckgiu6 = (Ozeiu6 & Azeiu6);
assign Azeiu6 = (Mwgiu6 & Twgiu6);
assign Twgiu6 = (Axgiu6 & Hxgiu6);
assign Hxgiu6 = (Oxgiu6 & Vxgiu6);
assign Vxgiu6 = (~(Cygiu6 | Tzfpw6[7]));
assign Cygiu6 = (Tzfpw6[8] | Tzfpw6[9]);
assign Oxgiu6 = (~(Jygiu6 | Tzfpw6[4]));
assign Jygiu6 = (Tzfpw6[5] | Tzfpw6[6]);
assign Axgiu6 = (Qygiu6 & Xygiu6);
assign Xygiu6 = (~(Ezgiu6 | Tzfpw6[23]));
assign Ezgiu6 = (Tzfpw6[2] | Tzfpw6[3]);
assign Qygiu6 = (~(Lzgiu6 | Tzfpw6[20]));
assign Lzgiu6 = (Tzfpw6[21] | Tzfpw6[22]);
assign Mwgiu6 = (Szgiu6 & Zzgiu6);
assign Zzgiu6 = (G0hiu6 & N0hiu6);
assign N0hiu6 = (~(U0hiu6 | Tzfpw6[18]));
assign U0hiu6 = (Tzfpw6[19] | Tzfpw6[1]);
assign G0hiu6 = (~(B1hiu6 | Tzfpw6[15]));
assign B1hiu6 = (Tzfpw6[16] | Tzfpw6[17]);
assign Szgiu6 = (I1hiu6 & P1hiu6);
assign P1hiu6 = (~(W1hiu6 | Tzfpw6[12]));
assign W1hiu6 = (Tzfpw6[13] | Tzfpw6[14]);
assign I1hiu6 = (~(Tzfpw6[10] | Tzfpw6[11]));
assign Ozeiu6 = (D2hiu6 & Bxghu6);
assign D2hiu6 = (Gc5iu6 & K2hiu6);
assign K2hiu6 = (R2hiu6 | STCALIB[25]);
assign R2hiu6 = (Ftghu6 | STCLKEN);
assign Djthu6 = (~(Y2hiu6 & F3hiu6));
assign F3hiu6 = (M3hiu6 & T3hiu6);
assign T3hiu6 = (~(HRDATA[7] & Pp7iu6));
assign M3hiu6 = (A4hiu6 & H4hiu6);
assign H4hiu6 = (~(Hrfpw6[7] & Uy4iu6));
assign A4hiu6 = (~(HRDATA[23] & Kq7iu6));
assign Y2hiu6 = (O4hiu6 & V4hiu6);
assign V4hiu6 = (~(Fr7iu6 & Df4iu6));
assign O4hiu6 = (C5hiu6 & J5hiu6);
assign J5hiu6 = (~(A25iu6 & Ppfpw6[7]));
assign C5hiu6 = (~(R05iu6 & D7fpw6[7]));
assign Withu6 = (~(Q5hiu6 & X5hiu6));
assign X5hiu6 = (E6hiu6 & L6hiu6);
assign L6hiu6 = (~(HRDATA[6] & Pp7iu6));
assign E6hiu6 = (S6hiu6 & Z6hiu6);
assign Z6hiu6 = (~(Hrfpw6[6] & Uy4iu6));
assign S6hiu6 = (~(HRDATA[22] & Kq7iu6));
assign Q5hiu6 = (G7hiu6 & N7hiu6);
assign N7hiu6 = (~(A25iu6 & Ppfpw6[6]));
assign G7hiu6 = (~(R05iu6 & D7fpw6[6]));
assign Pithu6 = (~(U7hiu6 & B8hiu6));
assign B8hiu6 = (I8hiu6 & P8hiu6);
assign P8hiu6 = (~(HRDATA[5] & Pp7iu6));
assign I8hiu6 = (W8hiu6 & D9hiu6);
assign D9hiu6 = (~(Hrfpw6[5] & Uy4iu6));
assign W8hiu6 = (~(HRDATA[21] & Kq7iu6));
assign U7hiu6 = (K9hiu6 & R9hiu6);
assign R9hiu6 = (~(Ppfpw6[5] & A25iu6));
assign K9hiu6 = (~(R05iu6 & D7fpw6[5]));
assign Iithu6 = (~(Y9hiu6 & Fahiu6));
assign Fahiu6 = (Mahiu6 & Tahiu6);
assign Tahiu6 = (~(HRDATA[4] & Pp7iu6));
assign Mahiu6 = (Abhiu6 & Hbhiu6);
assign Hbhiu6 = (~(Hrfpw6[4] & Uy4iu6));
assign Abhiu6 = (~(HRDATA[20] & Kq7iu6));
assign Y9hiu6 = (Obhiu6 & Vbhiu6);
assign Vbhiu6 = (~(Ppfpw6[4] & A25iu6));
assign Obhiu6 = (~(R05iu6 & D7fpw6[4]));
assign Bithu6 = (~(Cchiu6 & Jchiu6));
assign Jchiu6 = (Qchiu6 & Xchiu6);
assign Xchiu6 = (~(HRDATA[3] & Pp7iu6));
assign Qchiu6 = (Edhiu6 & Ldhiu6);
assign Ldhiu6 = (~(Hrfpw6[3] & Uy4iu6));
assign Edhiu6 = (~(HRDATA[19] & Kq7iu6));
assign Cchiu6 = (Sdhiu6 & Zdhiu6);
assign Zdhiu6 = (~(Fr7iu6 & H34iu6));
assign Sdhiu6 = (Gehiu6 & Nehiu6);
assign Nehiu6 = (~(Ppfpw6[3] & A25iu6));
assign Gehiu6 = (~(R05iu6 & D7fpw6[3]));
assign Uhthu6 = (~(Uehiu6 & Bfhiu6));
assign Bfhiu6 = (Ifhiu6 & Pfhiu6);
assign Pfhiu6 = (~(HRDATA[2] & Pp7iu6));
assign Ifhiu6 = (Wfhiu6 & Dghiu6);
assign Dghiu6 = (~(Hrfpw6[2] & Uy4iu6));
assign Wfhiu6 = (~(HRDATA[18] & Kq7iu6));
assign Uehiu6 = (Kghiu6 & Rghiu6);
assign Rghiu6 = (~(Fr7iu6 & Ud4iu6));
assign Kghiu6 = (Yghiu6 & Fhhiu6);
assign Fhhiu6 = (~(Ppfpw6[2] & A25iu6));
assign Yghiu6 = (~(R05iu6 & D7fpw6[2]));
assign Nhthu6 = (~(Mhhiu6 & Thhiu6));
assign Thhiu6 = (Aihiu6 & Hihiu6);
assign Hihiu6 = (~(HRDATA[1] & Pp7iu6));
assign Pp7iu6 = (Go7iu6 & M15iu6);
assign M15iu6 = (Oihiu6 & Vihiu6);
assign Oihiu6 = (Dxfhu6 & Cjhiu6);
assign Cjhiu6 = (~(vis_pc_o[0] & Jjhiu6));
assign Go7iu6 = (!T15iu6);
assign Aihiu6 = (Qjhiu6 & Xjhiu6);
assign Xjhiu6 = (~(Hrfpw6[1] & Uy4iu6));
assign Uy4iu6 = (Ekhiu6 & Vihiu6);
assign Ekhiu6 = (~(Lkhiu6 | Dxfhu6));
assign Lkhiu6 = (Pkciu6 & Skhiu6);
assign Skhiu6 = (Zkhiu6 | Ntfhu6);
assign Qjhiu6 = (~(HRDATA[17] & Kq7iu6));
assign Kq7iu6 = (Glhiu6 & Pz4iu6);
assign Pz4iu6 = (Nlhiu6 & Vihiu6);
assign Nlhiu6 = (vis_pc_o[0] & Jjhiu6);
assign Mhhiu6 = (Ulhiu6 & Bmhiu6);
assign Bmhiu6 = (Iz4iu6 | A34iu6);
assign Ulhiu6 = (Imhiu6 & Pmhiu6);
assign Pmhiu6 = (~(Ppfpw6[1] & A25iu6));
assign A25iu6 = (Ntfhu6 & Vihiu6);
assign Vihiu6 = (~(Wofiu6 | R05iu6));
assign Imhiu6 = (~(R05iu6 & D7fpw6[1]));
assign R05iu6 = (Wmhiu6 & Iz4iu6);
assign Iz4iu6 = (!Fr7iu6);
assign Fr7iu6 = (Dnhiu6 & Knhiu6);
assign Knhiu6 = (Rnhiu6 & Ynhiu6);
assign Rnhiu6 = (~(Jkgiu6 | Jfgpw6[4]));
assign Jkgiu6 = (!Npdhu6);
assign Dnhiu6 = (HALTED & Rzciu6);
assign Wmhiu6 = (~(Fohiu6 & Mohiu6));
assign Mohiu6 = (Tohiu6 & Aphiu6);
assign Tohiu6 = (Hphiu6 & Ophiu6);
assign Hphiu6 = (~(Vphiu6 & Cqhiu6));
assign Cqhiu6 = (Jqhiu6 | Qqhiu6);
assign Jqhiu6 = (~(Pkciu6 & Juzhu6));
assign Vphiu6 = (Eh6iu6 | Jjhiu6);
assign Fohiu6 = (Xqhiu6 & Erhiu6);
assign Xqhiu6 = (Lrhiu6 & Srhiu6);
assign Ghthu6 = (~(Zrhiu6 & Gshiu6));
assign Gshiu6 = (~(Nshiu6 & R6hhu6));
assign Nshiu6 = (Xbbiu6 & Jbbiu6);
assign Jbbiu6 = (!Mu4iu6);
assign Mu4iu6 = (Ushiu6 & Bthiu6);
assign Bthiu6 = (Ithiu6 & Pthiu6);
assign Ithiu6 = (~(Cyfpw6[7] | H4ghu6));
assign Ushiu6 = (~(Wthiu6 | Qjaiu6));
assign Xbbiu6 = (Duhiu6 | A2nhu6);
assign Zgthu6 = (Kuhiu6 & Ruhiu6);
assign Ruhiu6 = (Yuhiu6 & Fvhiu6);
assign Yuhiu6 = (~(Atdpw6 & Mvhiu6));
assign Kuhiu6 = (IRQ[16] & Tvhiu6);
assign Tvhiu6 = (~(Tk7iu6 & Awhiu6));
assign Awhiu6 = (Hwhiu6 | Qg6iu6);
assign Sgthu6 = (Owhiu6 & Vwhiu6);
assign Vwhiu6 = (Cxhiu6 & Jxhiu6);
assign Cxhiu6 = (~(Zvdpw6 & Qxhiu6));
assign Owhiu6 = (IRQ[30] & Xxhiu6);
assign Xxhiu6 = (~(Tk7iu6 & Eyhiu6));
assign Eyhiu6 = (Lyhiu6 | Qg6iu6);
assign Qg6iu6 = (!Fjfiu6);
assign Tk7iu6 = (~(Uc5iu6 & Fjfiu6));
assign Fjfiu6 = (~(Syhiu6 & Zyhiu6));
assign Zyhiu6 = (Gzhiu6 & Nzhiu6);
assign Gzhiu6 = (~(Ur4iu6 | Gc5iu6));
assign Syhiu6 = (I4eiu6 & Uzhiu6);
assign Lgthu6 = (~(B0iiu6 & I0iiu6));
assign I0iiu6 = (P0iiu6 & W0iiu6);
assign W0iiu6 = (~(vis_pc_o[3] & Ok8iu6));
assign P0iiu6 = (D1iiu6 & K1iiu6);
assign K1iiu6 = (~(Jl8iu6 & Tugpw6[2]));
assign Tugpw6[2] = (~(R1iiu6 & Y1iiu6));
assign Y1iiu6 = (~(N5fpw6[3] & Sdaiu6));
assign R1iiu6 = (F2iiu6 & M2iiu6);
assign M2iiu6 = (T2iiu6 | Eg0iu6);
assign F2iiu6 = (~(Eafpw6[4] & A3iiu6));
assign D1iiu6 = (~(Ql8iu6 & vis_ipsr_o[4]));
assign B0iiu6 = (H3iiu6 & O3iiu6);
assign O3iiu6 = (Lm8iu6 | V3iiu6);
assign H3iiu6 = (~(Zm8iu6 & H34iu6));
assign Egthu6 = (~(C4iiu6 & J4iiu6));
assign J4iiu6 = (Q4iiu6 & X4iiu6);
assign X4iiu6 = (~(Ok8iu6 & vis_pc_o[1]));
assign Q4iiu6 = (E5iiu6 & L5iiu6);
assign L5iiu6 = (~(Jl8iu6 & Tugpw6[0]));
assign Tugpw6[0] = (~(S5iiu6 & Z5iiu6));
assign Z5iiu6 = (~(Eafpw6[2] & A3iiu6));
assign S5iiu6 = (G6iiu6 & N6iiu6);
assign N6iiu6 = (~(Sdaiu6 & U6iiu6));
assign U6iiu6 = (Vtzhu6 ^ Cuzhu6);
assign Cuzhu6 = (Juzhu6 ^ Quzhu6);
assign G6iiu6 = (~(B7iiu6 & Gh0iu6));
assign E5iiu6 = (~(Ql8iu6 & vis_ipsr_o[2]));
assign C4iiu6 = (I7iiu6 & P7iiu6);
assign P7iiu6 = (~(W29iu6 & Fkfpw6[2]));
assign I7iiu6 = (~(Zm8iu6 & Ud4iu6));
assign Xfthu6 = (D8iiu6 ? W7iiu6 : S8fpw6[8]);
assign W7iiu6 = (~(K8iiu6 & R8iiu6));
assign R8iiu6 = (Y8iiu6 & F9iiu6);
assign F9iiu6 = (~(D7fpw6[0] & M9iiu6));
assign Y8iiu6 = (~(D7fpw6[8] & T9iiu6));
assign K8iiu6 = (Aaiiu6 & Haiiu6);
assign Haiiu6 = (Oaiiu6 | O95iu6);
assign Qfthu6 = (~(Vaiiu6 & Cbiiu6));
assign Cbiiu6 = (~(Jbiiu6 & Qbiiu6));
assign Vaiiu6 = (D8iiu6 ? Xbiiu6 : P65iu6);
assign Xbiiu6 = (Eciiu6 & Lciiu6);
assign Lciiu6 = (Sciiu6 & Zciiu6);
assign Zciiu6 = (~(D7fpw6[1] & M9iiu6));
assign Sciiu6 = (~(D7fpw6[9] & T9iiu6));
assign Eciiu6 = (Aaiiu6 & Gdiiu6);
assign Gdiiu6 = (Oaiiu6 | Ndiiu6);
assign Jfthu6 = (~(Udiiu6 & Beiiu6));
assign Beiiu6 = (~(S8fpw6[10] & Ieiiu6));
assign Ieiiu6 = (~(D8iiu6 & Peiiu6));
assign Peiiu6 = (~(Jbiiu6 & Weiiu6));
assign Jbiiu6 = (~(Dfiiu6 | Kfiiu6));
assign Udiiu6 = (~(D8iiu6 & Rfiiu6));
assign Rfiiu6 = (~(Yfiiu6 & Fgiiu6));
assign Fgiiu6 = (Mgiiu6 & Tgiiu6);
assign Tgiiu6 = (~(D7fpw6[2] & M9iiu6));
assign M9iiu6 = (~(Ahiiu6 & Hhiiu6));
assign Hhiiu6 = (Ohiiu6 & Vhiiu6);
assign Ohiiu6 = (~(Ciiiu6 & Jiiiu6));
assign Ciiiu6 = (Qiiiu6 & Zraiu6);
assign Qiiiu6 = (Xiiiu6 | Ejiiu6);
assign Ahiiu6 = (Ljiiu6 & Sjiiu6);
assign Sjiiu6 = (Zjiiu6 | Gkiiu6);
assign Mgiiu6 = (~(D7fpw6[10] & T9iiu6));
assign T9iiu6 = (~(Nkiiu6 & Ukiiu6));
assign Ukiiu6 = (Bliiu6 & Iliiu6);
assign Iliiu6 = (~(Pliiu6 & Wliiu6));
assign Pliiu6 = (Dmiiu6 & Zraiu6);
assign Bliiu6 = (~(Kmiiu6 | Rmiiu6));
assign Nkiiu6 = (Ymiiu6 & Fniiu6);
assign Yfiiu6 = (Aaiiu6 & Mniiu6);
assign Mniiu6 = (Oaiiu6 | Tniiu6);
assign Cfthu6 = (Aoiiu6 | Hoiiu6);
assign Hoiiu6 = (~(Ooiiu6 | Voiiu6));
assign Ooiiu6 = (Dfiiu6 | Kfiiu6);
assign Dfiiu6 = (~(Y7ghu6 | U98iu6));
assign Aoiiu6 = (D8iiu6 ? Cpiiu6 : S8fpw6[11]);
assign D8iiu6 = (HREADY & Jpiiu6);
assign Jpiiu6 = (~(Qpiiu6 & Xpiiu6));
assign Xpiiu6 = (Eqiiu6 & Lqiiu6);
assign Lqiiu6 = (Sqiiu6 & Zqiiu6);
assign Zqiiu6 = (~(Griiu6 & Nriiu6));
assign Griiu6 = (~(Uriiu6 | Y7ghu6));
assign Sqiiu6 = (Bsiiu6 & Isiiu6);
assign Bsiiu6 = (~(Psiiu6 & Ae0iu6));
assign Psiiu6 = (~(Mjfiu6 | H4ghu6));
assign Eqiiu6 = (Wsiiu6 & Dtiiu6);
assign Dtiiu6 = (~(Ktiiu6 & Ndiiu6));
assign Ktiiu6 = (~(Rtiiu6 & Ytiiu6));
assign Ytiiu6 = (~(D7fpw6[10] & Fuiiu6));
assign Fuiiu6 = (~(Muiiu6 & Tuiiu6));
assign Tuiiu6 = (~(Aviiu6 & Hviiu6));
assign Aviiu6 = (~(Oviiu6 | Zwciu6));
assign Muiiu6 = (~(Vviiu6 & Cwiiu6));
assign Rtiiu6 = (~(Vviiu6 & Jwiiu6));
assign Wsiiu6 = (Qwiiu6 & Xwiiu6);
assign Xwiiu6 = (~(D7fpw6[14] & Exiiu6));
assign Exiiu6 = (~(Lxiiu6 & Sxiiu6));
assign Sxiiu6 = (~(Zxiiu6 & C0ehu6));
assign Zxiiu6 = (Gyiiu6 & Q5aiu6);
assign Gyiiu6 = (S1ehu6 | Nyiiu6);
assign Lxiiu6 = (~(Ejiiu6 & Uyiiu6));
assign Qwiiu6 = (~(Bziiu6 & Uyiiu6));
assign Qpiiu6 = (Iziiu6 & Pziiu6);
assign Pziiu6 = (Wziiu6 & D0jiu6);
assign Wziiu6 = (K0jiu6 & R0jiu6);
assign R0jiu6 = (~(Y0jiu6 & F1jiu6));
assign Iziiu6 = (M1jiu6 & T1jiu6);
assign Cpiiu6 = (~(A2jiu6 & H2jiu6));
assign H2jiu6 = (O2jiu6 & V2jiu6);
assign V2jiu6 = (~(D7fpw6[11] & C3jiu6));
assign C3jiu6 = (Kmiiu6 | J3jiu6);
assign J3jiu6 = (Rmiiu6 & D7fpw6[12]);
assign Kmiiu6 = (Zraiu6 & Q3jiu6);
assign Q3jiu6 = (~(X3jiu6 & E4jiu6));
assign O2jiu6 = (V4aiu6 | Ljiiu6);
assign Ljiiu6 = (L4jiu6 & S4jiu6);
assign L4jiu6 = (~(Z4jiu6 & G5jiu6));
assign G5jiu6 = (N5jiu6 & U5jiu6);
assign N5jiu6 = (Oviiu6 | Tniiu6);
assign A2jiu6 = (Aaiiu6 & B6jiu6);
assign B6jiu6 = (Oaiiu6 | I6jiu6);
assign Aaiiu6 = (P6jiu6 & W6jiu6);
assign P6jiu6 = (D7jiu6 & Faaiu6);
assign D7jiu6 = (~(K7jiu6 & R7jiu6));
assign K7jiu6 = (Ia8iu6 & D7fpw6[7]);
assign Vethu6 = (F58iu6 ? S8fpw6[3] : Y7jiu6);
assign Y7jiu6 = (~(F8jiu6 & M8jiu6));
assign M8jiu6 = (T8jiu6 & A9jiu6);
assign A9jiu6 = (H9jiu6 & O9jiu6);
assign O9jiu6 = (~(V9jiu6 & Ce8iu6));
assign V9jiu6 = (~(Cajiu6 ^ Jajiu6));
assign Jajiu6 = (Qajiu6 & S8fpw6[2]);
assign H9jiu6 = (Xajiu6 & Faaiu6);
assign Xajiu6 = (~(Ebjiu6 & E88iu6));
assign Ebjiu6 = (~(Lbjiu6 & Sbjiu6));
assign Sbjiu6 = (~(Zbjiu6 & Gcjiu6));
assign Lbjiu6 = (~(Ncjiu6 & Ucjiu6));
assign T8jiu6 = (Bdjiu6 & Idjiu6);
assign Idjiu6 = (~(Tc8iu6 & Ppfpw6[3]));
assign Bdjiu6 = (~(D7fpw6[9] & Pdjiu6));
assign F8jiu6 = (Wdjiu6 & Dejiu6);
assign Dejiu6 = (Kejiu6 & Rejiu6);
assign Rejiu6 = (~(Habiu6 & D7fpw6[2]));
assign Kejiu6 = (V4aiu6 | Yb8iu6);
assign Wdjiu6 = (Yejiu6 & Ffjiu6);
assign Ffjiu6 = (~(Cbbiu6 & D7fpw6[8]));
assign Yejiu6 = (~(Mfjiu6 & Tfjiu6));
assign Oethu6 = (F58iu6 ? S8fpw6[2] : Agjiu6);
assign F58iu6 = (~(HREADY & Hgjiu6));
assign Hgjiu6 = (~(Ogjiu6 & Vgjiu6));
assign Vgjiu6 = (Chjiu6 & Jhjiu6);
assign Jhjiu6 = (Qhjiu6 & Xhjiu6);
assign Xhjiu6 = (~(Eijiu6 & Lijiu6));
assign Eijiu6 = (~(Sijiu6 | Cyfpw6[0]));
assign Qhjiu6 = (Zijiu6 & Gjjiu6);
assign Zijiu6 = (~(Njjiu6 & Ujjiu6));
assign Njjiu6 = (~(Q5aiu6 | Bkjiu6));
assign Chjiu6 = (Ikjiu6 & Pkjiu6);
assign Pkjiu6 = (~(Wkjiu6 & D7fpw6[10]));
assign Ikjiu6 = (Dljiu6 & Kljiu6);
assign Kljiu6 = (~(Rljiu6 & Yljiu6));
assign Dljiu6 = (Fmjiu6 | Mmjiu6);
assign Ogjiu6 = (Tmjiu6 & Anjiu6);
assign Anjiu6 = (Hnjiu6 & Onjiu6);
assign Hnjiu6 = (Vnjiu6 & Cojiu6);
assign Cojiu6 = (Wmaiu6 | Jojiu6);
assign Vnjiu6 = (Qojiu6 | Xojiu6);
assign Tmjiu6 = (Epjiu6 & Lpjiu6);
assign Lpjiu6 = (~(Ae0iu6 & Pthiu6));
assign Agjiu6 = (~(Spjiu6 & Zpjiu6));
assign Zpjiu6 = (Gqjiu6 & Nqjiu6);
assign Nqjiu6 = (Uqjiu6 & V68iu6);
assign V68iu6 = (~(W8aiu6 & Brjiu6));
assign Brjiu6 = (~(Irjiu6 & Wthiu6));
assign Irjiu6 = (Prjiu6 | Cyfpw6[5]);
assign Uqjiu6 = (~(Wrjiu6 & E88iu6));
assign E88iu6 = (~(Dsjiu6 & Ksjiu6));
assign Ksjiu6 = (~(Rsjiu6 & Ysjiu6));
assign Ysjiu6 = (~(Oviiu6 | Ftjiu6));
assign Rsjiu6 = (Ia8iu6 & Mtjiu6);
assign Dsjiu6 = (~(Ttjiu6 & Aujiu6));
assign Ttjiu6 = (~(Hujiu6 | I6jiu6));
assign Wrjiu6 = (Gcjiu6 ^ Zbjiu6);
assign Zbjiu6 = (W7biu6 & P7biu6);
assign P7biu6 = (~(Oujiu6 | Ncjiu6));
assign Oujiu6 = (Vujiu6 & Cvjiu6);
assign W7biu6 = (L88iu6 & S88iu6);
assign S88iu6 = (Jvjiu6 ^ O95iu6);
assign Gcjiu6 = (Ucjiu6 ^ Ncjiu6);
assign Ncjiu6 = (~(Cvjiu6 | Vujiu6));
assign Vujiu6 = (~(Qvjiu6 & Xvjiu6));
assign Xvjiu6 = (Ewjiu6 | Lwjiu6);
assign Cvjiu6 = (O95iu6 | Jvjiu6);
assign Jvjiu6 = (Swjiu6 ^ D7fpw6[6]);
assign Ucjiu6 = (~(Zwjiu6 & Gxjiu6));
assign Gxjiu6 = (Nxjiu6 & Qvjiu6);
assign Qvjiu6 = (~(Lwjiu6 & Ewjiu6));
assign Ewjiu6 = (Uxjiu6 ^ Byjiu6);
assign Lwjiu6 = (~(Ad8iu6 | Swjiu6));
assign Swjiu6 = (Iyjiu6 ^ D7fpw6[5]);
assign Nxjiu6 = (~(Byjiu6 & Uxjiu6));
assign Uxjiu6 = (Pyjiu6 ^ Wyjiu6);
assign Byjiu6 = (~(Dzjiu6 | Iyjiu6));
assign Iyjiu6 = (Kzjiu6 ^ D7fpw6[4]);
assign Zwjiu6 = (Rzjiu6 & Yzjiu6);
assign Yzjiu6 = (~(Wyjiu6 & Pyjiu6));
assign Pyjiu6 = (~(F0kiu6 ^ M0kiu6));
assign F0kiu6 = (V4aiu6 | T0kiu6);
assign Wyjiu6 = (~(A1kiu6 | Kzjiu6));
assign Kzjiu6 = (H1kiu6 ^ V4aiu6);
assign Rzjiu6 = (~(O1kiu6 & D7fpw6[3]));
assign O1kiu6 = (H1kiu6 & M0kiu6);
assign M0kiu6 = (~(V1kiu6 & C2kiu6));
assign C2kiu6 = (Prjiu6 | J2kiu6);
assign V1kiu6 = (Rb8iu6 | Ccaiu6);
assign H1kiu6 = (!T0kiu6);
assign T0kiu6 = (J2kiu6 ^ D7fpw6[2]);
assign J2kiu6 = (~(D7fpw6[0] ^ D7fpw6[1]));
assign Gqjiu6 = (Q2kiu6 & X2kiu6);
assign X2kiu6 = (~(E3kiu6 & Ce8iu6));
assign Ce8iu6 = (~(L3kiu6 & S3kiu6));
assign L3kiu6 = (Z3kiu6 & G4kiu6);
assign G4kiu6 = (~(N4kiu6 & Cyfpw6[5]));
assign Z3kiu6 = (~(U98iu6 & U4kiu6));
assign E3kiu6 = (~(B5kiu6 ^ Qajiu6));
assign Qajiu6 = (~(Je8iu6 | Y8biu6));
assign Q2kiu6 = (~(Tc8iu6 & Ppfpw6[2]));
assign Tc8iu6 = (Ivfhu6 & I5kiu6);
assign I5kiu6 = (~(P5kiu6 & W5kiu6));
assign W5kiu6 = (~(D6kiu6 & Qjaiu6));
assign Spjiu6 = (K6kiu6 & R6kiu6);
assign R6kiu6 = (Y6kiu6 & F7kiu6);
assign F7kiu6 = (Ndiiu6 | Hd8iu6);
assign Hd8iu6 = (~(Pdjiu6 | M7kiu6));
assign Pdjiu6 = (~(T7kiu6 & A8kiu6));
assign A8kiu6 = (~(H8kiu6 & Ftjiu6));
assign H8kiu6 = (~(O8kiu6 & Vhiiu6));
assign T7kiu6 = (~(M7kiu6 & Oviiu6));
assign Y6kiu6 = (~(Habiu6 & D7fpw6[1]));
assign Habiu6 = (Ia8iu6 & V8kiu6);
assign V8kiu6 = (~(H95iu6 & C9kiu6));
assign C9kiu6 = (~(J9kiu6 & Oviiu6));
assign K6kiu6 = (Q9kiu6 & X9kiu6);
assign X9kiu6 = (Prjiu6 | Yb8iu6);
assign Yb8iu6 = (Eakiu6 & Lakiu6);
assign Lakiu6 = (Sakiu6 & Zjiiu6);
assign Zjiiu6 = (!Zakiu6);
assign Sakiu6 = (~(Gbkiu6 & Nyiiu6));
assign Gbkiu6 = (Ia8iu6 & Nbkiu6);
assign Eakiu6 = (Ubkiu6 & Bckiu6);
assign Bckiu6 = (E4jiu6 | Jcaiu6);
assign Q9kiu6 = (~(Cbbiu6 & D7fpw6[7]));
assign Hethu6 = (Ickiu6 ? vis_r2_o[2] : Qcaiu6);
assign Aethu6 = (Ickiu6 ? vis_r2_o[4] : Ef8iu6);
assign Tdthu6 = (Ickiu6 ? vis_r2_o[23] : Vx9iu6);
assign Mdthu6 = (Ickiu6 ? vis_r2_o[30] : K39iu6);
assign Fdthu6 = (Ickiu6 ? vis_r2_o[31] : D39iu6);
assign Ycthu6 = (Ickiu6 ? vis_r2_o[0] : Tx8iu6);
assign Rcthu6 = (Pckiu6 ? vis_r3_o[2] : Qcaiu6);
assign Kcthu6 = (Pckiu6 ? vis_r3_o[4] : Ef8iu6);
assign Dcthu6 = (Pckiu6 ? vis_r3_o[23] : Vx9iu6);
assign Wbthu6 = (Pckiu6 ? vis_r3_o[30] : K39iu6);
assign Pbthu6 = (Pckiu6 ? vis_r3_o[31] : D39iu6);
assign Ibthu6 = (Pckiu6 ? vis_r3_o[0] : Tx8iu6);
assign Bbthu6 = (Wckiu6 ? vis_r4_o[2] : Qcaiu6);
assign Uathu6 = (Wckiu6 ? vis_r4_o[4] : Ef8iu6);
assign Nathu6 = (Wckiu6 ? vis_r4_o[23] : Vx9iu6);
assign Gathu6 = (Wckiu6 ? vis_r4_o[30] : K39iu6);
assign Z9thu6 = (Wckiu6 ? vis_r4_o[31] : D39iu6);
assign S9thu6 = (Wckiu6 ? vis_r4_o[0] : Tx8iu6);
assign L9thu6 = (Ddkiu6 ? vis_r5_o[2] : Qcaiu6);
assign E9thu6 = (Ddkiu6 ? vis_r5_o[4] : Ef8iu6);
assign X8thu6 = (Ddkiu6 ? vis_r5_o[23] : Vx9iu6);
assign Q8thu6 = (Ddkiu6 ? vis_r5_o[30] : K39iu6);
assign J8thu6 = (Ddkiu6 ? vis_r5_o[31] : D39iu6);
assign C8thu6 = (Ddkiu6 ? vis_r5_o[0] : Tx8iu6);
assign V7thu6 = (Kdkiu6 ? vis_r6_o[2] : Qcaiu6);
assign O7thu6 = (Kdkiu6 ? vis_r6_o[4] : Ef8iu6);
assign H7thu6 = (Kdkiu6 ? vis_r6_o[23] : Vx9iu6);
assign A7thu6 = (Kdkiu6 ? vis_r6_o[30] : K39iu6);
assign T6thu6 = (Kdkiu6 ? vis_r6_o[31] : D39iu6);
assign M6thu6 = (Kdkiu6 ? vis_r6_o[0] : Tx8iu6);
assign F6thu6 = (Rdkiu6 ? vis_r7_o[2] : Qcaiu6);
assign Y5thu6 = (Rdkiu6 ? vis_r7_o[4] : Ef8iu6);
assign R5thu6 = (Rdkiu6 ? vis_r7_o[23] : Vx9iu6);
assign K5thu6 = (Rdkiu6 ? vis_r7_o[30] : K39iu6);
assign D5thu6 = (Rdkiu6 ? vis_r7_o[31] : D39iu6);
assign W4thu6 = (Rdkiu6 ? vis_r7_o[0] : Tx8iu6);
assign P4thu6 = (Ydkiu6 ? Qcaiu6 : vis_psp_o[0]);
assign I4thu6 = (Ydkiu6 ? D39iu6 : vis_psp_o[29]);
assign B4thu6 = (Ydkiu6 ? K39iu6 : vis_psp_o[28]);
assign U3thu6 = (Ydkiu6 ? Vx9iu6 : vis_psp_o[21]);
assign N3thu6 = (Ydkiu6 ? Ef8iu6 : vis_psp_o[2]);
assign G3thu6 = (Fekiu6 ? Qcaiu6 : vis_msp_o[0]);
assign Z2thu6 = (Fekiu6 ? D39iu6 : vis_msp_o[29]);
assign S2thu6 = (Fekiu6 ? K39iu6 : vis_msp_o[28]);
assign L2thu6 = (Fekiu6 ? Vx9iu6 : vis_msp_o[21]);
assign E2thu6 = (Fekiu6 ? Ef8iu6 : vis_msp_o[2]);
assign X1thu6 = (Mekiu6 ? vis_r14_o[2] : Qcaiu6);
assign Q1thu6 = (Mekiu6 ? vis_r14_o[4] : Ef8iu6);
assign J1thu6 = (Mekiu6 ? vis_r14_o[23] : Vx9iu6);
assign C1thu6 = (Mekiu6 ? vis_r14_o[30] : K39iu6);
assign V0thu6 = (Mekiu6 ? vis_r14_o[31] : D39iu6);
assign O0thu6 = (Mekiu6 ? vis_r14_o[0] : Tx8iu6);
assign H0thu6 = (Tekiu6 ? vis_r12_o[2] : Qcaiu6);
assign A0thu6 = (Tekiu6 ? vis_r12_o[4] : Ef8iu6);
assign Tzshu6 = (Tekiu6 ? vis_r12_o[23] : Vx9iu6);
assign Mzshu6 = (Tekiu6 ? vis_r12_o[30] : K39iu6);
assign Fzshu6 = (Tekiu6 ? vis_r12_o[31] : D39iu6);
assign Yyshu6 = (Tekiu6 ? vis_r12_o[0] : Tx8iu6);
assign Ryshu6 = (Afkiu6 ? vis_r11_o[2] : Qcaiu6);
assign Kyshu6 = (Afkiu6 ? vis_r11_o[4] : Ef8iu6);
assign Dyshu6 = (Afkiu6 ? vis_r11_o[23] : Vx9iu6);
assign Wxshu6 = (Afkiu6 ? vis_r11_o[30] : K39iu6);
assign Pxshu6 = (Afkiu6 ? vis_r11_o[31] : D39iu6);
assign Ixshu6 = (Afkiu6 ? vis_r11_o[0] : Tx8iu6);
assign Bxshu6 = (Hfkiu6 ? vis_r10_o[2] : Qcaiu6);
assign Uwshu6 = (Hfkiu6 ? vis_r10_o[4] : Ef8iu6);
assign Nwshu6 = (Hfkiu6 ? vis_r10_o[23] : Vx9iu6);
assign Gwshu6 = (Hfkiu6 ? vis_r10_o[30] : K39iu6);
assign Zvshu6 = (Hfkiu6 ? vis_r10_o[31] : D39iu6);
assign Svshu6 = (Hfkiu6 ? vis_r10_o[0] : Tx8iu6);
assign Lvshu6 = (Ofkiu6 ? vis_r9_o[2] : Qcaiu6);
assign Evshu6 = (Ofkiu6 ? vis_r9_o[4] : Ef8iu6);
assign Xushu6 = (Ofkiu6 ? vis_r9_o[23] : Vx9iu6);
assign Qushu6 = (Ofkiu6 ? vis_r9_o[30] : K39iu6);
assign Jushu6 = (Ofkiu6 ? vis_r9_o[31] : D39iu6);
assign Cushu6 = (Ofkiu6 ? vis_r9_o[0] : Tx8iu6);
assign Vtshu6 = (Vfkiu6 ? vis_r8_o[2] : Qcaiu6);
assign Qcaiu6 = (~(Ogciu6 & Cgkiu6));
assign Otshu6 = (Vfkiu6 ? vis_r8_o[3] : Jgkiu6);
assign Htshu6 = (~(Qgkiu6 & Xgkiu6));
assign Xgkiu6 = (Ehkiu6 & Lhkiu6);
assign Lhkiu6 = (~(Ok8iu6 & vis_pc_o[2]));
assign Ehkiu6 = (Shkiu6 & Zhkiu6);
assign Zhkiu6 = (~(Jl8iu6 & Tugpw6[1]));
assign Tugpw6[1] = (~(Gikiu6 & Nikiu6));
assign Nikiu6 = (~(N5fpw6[2] & Sdaiu6));
assign Gikiu6 = (Uikiu6 & Bjkiu6);
assign Bjkiu6 = (T2iiu6 | Lg0iu6);
assign Uikiu6 = (~(Eafpw6[3] & A3iiu6));
assign Shkiu6 = (~(Ql8iu6 & vis_ipsr_o[3]));
assign Qgkiu6 = (Ijkiu6 & Pjkiu6);
assign Pjkiu6 = (Lm8iu6 | Wjkiu6);
assign Ijkiu6 = (~(Zm8iu6 & Df4iu6));
assign Atshu6 = (Ydkiu6 ? Jgkiu6 : vis_psp_o[1]);
assign Tsshu6 = (Fekiu6 ? Jgkiu6 : vis_msp_o[1]);
assign Msshu6 = (Mekiu6 ? vis_r14_o[3] : Jgkiu6);
assign Fsshu6 = (Tekiu6 ? vis_r12_o[3] : Jgkiu6);
assign Yrshu6 = (Rdkiu6 ? vis_r7_o[3] : Jgkiu6);
assign Rrshu6 = (Kdkiu6 ? vis_r6_o[3] : Jgkiu6);
assign Krshu6 = (Ddkiu6 ? vis_r5_o[3] : Jgkiu6);
assign Drshu6 = (Wckiu6 ? vis_r4_o[3] : Jgkiu6);
assign Wqshu6 = (Afkiu6 ? vis_r11_o[3] : Jgkiu6);
assign Pqshu6 = (Hfkiu6 ? vis_r10_o[3] : Jgkiu6);
assign Iqshu6 = (Ofkiu6 ? vis_r9_o[3] : Jgkiu6);
assign Bqshu6 = (Pckiu6 ? vis_r3_o[3] : Jgkiu6);
assign Upshu6 = (Ickiu6 ? vis_r2_o[3] : Jgkiu6);
assign Npshu6 = (Mx8iu6 ? vis_r1_o[3] : Jgkiu6);
assign Gpshu6 = (Lf8iu6 ? vis_r0_o[3] : Jgkiu6);
assign Jgkiu6 = (~(Kifiu6 & Dkkiu6));
assign Zoshu6 = (Vfkiu6 ? vis_r8_o[4] : Ef8iu6);
assign Ef8iu6 = (~(Y4fiu6 & Kkkiu6));
assign Soshu6 = (Vfkiu6 ? vis_r8_o[5] : Rkkiu6);
assign Loshu6 = (~(Ykkiu6 & Flkiu6));
assign Flkiu6 = (Mlkiu6 & Tlkiu6);
assign Tlkiu6 = (~(vis_pc_o[4] & Ok8iu6));
assign Mlkiu6 = (Amkiu6 & Hmkiu6);
assign Hmkiu6 = (~(Jl8iu6 & Tugpw6[3]));
assign Tugpw6[3] = (~(Omkiu6 & Vmkiu6));
assign Vmkiu6 = (~(N5fpw6[4] & Sdaiu6));
assign Omkiu6 = (Cnkiu6 & Jnkiu6);
assign Jnkiu6 = (T2iiu6 | Xf0iu6);
assign Cnkiu6 = (~(Eafpw6[5] & A3iiu6));
assign Amkiu6 = (~(Ql8iu6 & vis_ipsr_o[5]));
assign Ykkiu6 = (Qnkiu6 & Xnkiu6);
assign Xnkiu6 = (Lm8iu6 | Eokiu6);
assign Qnkiu6 = (~(Zm8iu6 & Oh4iu6));
assign Eoshu6 = (Ydkiu6 ? Rkkiu6 : vis_psp_o[3]);
assign Xnshu6 = (Fekiu6 ? Rkkiu6 : vis_msp_o[3]);
assign Qnshu6 = (Mekiu6 ? vis_r14_o[5] : Rkkiu6);
assign Jnshu6 = (Tekiu6 ? vis_r12_o[5] : Rkkiu6);
assign Cnshu6 = (Rdkiu6 ? vis_r7_o[5] : Rkkiu6);
assign Vmshu6 = (Kdkiu6 ? vis_r6_o[5] : Rkkiu6);
assign Omshu6 = (Ddkiu6 ? vis_r5_o[5] : Rkkiu6);
assign Hmshu6 = (Wckiu6 ? vis_r4_o[5] : Rkkiu6);
assign Amshu6 = (Afkiu6 ? vis_r11_o[5] : Rkkiu6);
assign Tlshu6 = (Hfkiu6 ? vis_r10_o[5] : Rkkiu6);
assign Mlshu6 = (Ofkiu6 ? vis_r9_o[5] : Rkkiu6);
assign Flshu6 = (Pckiu6 ? vis_r3_o[5] : Rkkiu6);
assign Ykshu6 = (Ickiu6 ? vis_r2_o[5] : Rkkiu6);
assign Rkshu6 = (Mx8iu6 ? vis_r1_o[5] : Rkkiu6);
assign Kkshu6 = (Lf8iu6 ? vis_r0_o[5] : Rkkiu6);
assign Rkkiu6 = (~(Ljbiu6 & Lokiu6));
assign Dkshu6 = (Vfkiu6 ? vis_r8_o[6] : Sokiu6);
assign Wjshu6 = (~(Zokiu6 & Gpkiu6));
assign Gpkiu6 = (Npkiu6 & Upkiu6);
assign Upkiu6 = (~(Jl8iu6 & Tugpw6[4]));
assign Npkiu6 = (~(vis_pc_o[5] & Ok8iu6));
assign Zokiu6 = (Bqkiu6 & Iqkiu6);
assign Iqkiu6 = (~(W29iu6 & Fkfpw6[6]));
assign Bqkiu6 = (~(Zm8iu6 & Xi4iu6));
assign Pjshu6 = (Ydkiu6 ? Sokiu6 : vis_psp_o[4]);
assign Ijshu6 = (Fekiu6 ? Sokiu6 : vis_msp_o[4]);
assign Bjshu6 = (Mekiu6 ? vis_r14_o[6] : Sokiu6);
assign Uishu6 = (Tekiu6 ? vis_r12_o[6] : Sokiu6);
assign Nishu6 = (Rdkiu6 ? vis_r7_o[6] : Sokiu6);
assign Gishu6 = (Kdkiu6 ? vis_r6_o[6] : Sokiu6);
assign Zhshu6 = (Ddkiu6 ? vis_r5_o[6] : Sokiu6);
assign Shshu6 = (Wckiu6 ? vis_r4_o[6] : Sokiu6);
assign Lhshu6 = (Afkiu6 ? vis_r11_o[6] : Sokiu6);
assign Ehshu6 = (Hfkiu6 ? vis_r10_o[6] : Sokiu6);
assign Xgshu6 = (Ofkiu6 ? vis_r9_o[6] : Sokiu6);
assign Qgshu6 = (Pckiu6 ? vis_r3_o[6] : Sokiu6);
assign Jgshu6 = (Ickiu6 ? vis_r2_o[6] : Sokiu6);
assign Cgshu6 = (Mx8iu6 ? vis_r1_o[6] : Sokiu6);
assign Vfshu6 = (Lf8iu6 ? vis_r0_o[6] : Sokiu6);
assign Sokiu6 = (Pqkiu6 | Wqkiu6);
assign Ofshu6 = (Vfkiu6 ? vis_r8_o[7] : Drkiu6);
assign Hfshu6 = (~(Krkiu6 & Rrkiu6));
assign Rrkiu6 = (Yrkiu6 & Fskiu6);
assign Fskiu6 = (~(Jl8iu6 & Tugpw6[5]));
assign Tugpw6[5] = (~(Mskiu6 & Tskiu6));
assign Tskiu6 = (~(N5fpw6[6] & Sdaiu6));
assign Mskiu6 = (Atkiu6 & Htkiu6);
assign Htkiu6 = (T2iiu6 | Jf0iu6);
assign Atkiu6 = (~(Eafpw6[7] & A3iiu6));
assign Yrkiu6 = (~(vis_pc_o[6] & Ok8iu6));
assign Krkiu6 = (Otkiu6 & Vtkiu6);
assign Vtkiu6 = (Lm8iu6 | Cukiu6);
assign Otkiu6 = (~(Zm8iu6 & Gk4iu6));
assign Afshu6 = (Ydkiu6 ? Drkiu6 : vis_psp_o[5]);
assign Teshu6 = (Fekiu6 ? Drkiu6 : vis_msp_o[5]);
assign Meshu6 = (Mekiu6 ? vis_r14_o[7] : Drkiu6);
assign Feshu6 = (Tekiu6 ? vis_r12_o[7] : Drkiu6);
assign Ydshu6 = (Rdkiu6 ? vis_r7_o[7] : Drkiu6);
assign Rdshu6 = (Kdkiu6 ? vis_r6_o[7] : Drkiu6);
assign Kdshu6 = (Ddkiu6 ? vis_r5_o[7] : Drkiu6);
assign Ddshu6 = (Wckiu6 ? vis_r4_o[7] : Drkiu6);
assign Wcshu6 = (Afkiu6 ? vis_r11_o[7] : Drkiu6);
assign Pcshu6 = (Hfkiu6 ? vis_r10_o[7] : Drkiu6);
assign Icshu6 = (Ofkiu6 ? vis_r9_o[7] : Drkiu6);
assign Bcshu6 = (Pckiu6 ? vis_r3_o[7] : Drkiu6);
assign Ubshu6 = (Ickiu6 ? vis_r2_o[7] : Drkiu6);
assign Nbshu6 = (Mx8iu6 ? vis_r1_o[7] : Drkiu6);
assign Gbshu6 = (Lf8iu6 ? vis_r0_o[7] : Drkiu6);
assign Drkiu6 = (Jukiu6 | Qukiu6);
assign Zashu6 = (Vfkiu6 ? vis_r8_o[23] : Vx9iu6);
assign Vx9iu6 = (~(Xukiu6 & Evkiu6));
assign Xukiu6 = (Lvkiu6 & Svkiu6);
assign Sashu6 = (Vfkiu6 ? vis_r8_o[24] : Zvkiu6);
assign Lashu6 = (~(Gwkiu6 & Nwkiu6));
assign Nwkiu6 = (Uwkiu6 & Bxkiu6);
assign Bxkiu6 = (~(vis_pc_o[23] & Ok8iu6));
assign Uwkiu6 = (Ixkiu6 & Pxkiu6);
assign Pxkiu6 = (~(Jl8iu6 & Tzdpw6));
assign Ixkiu6 = (~(Ql8iu6 & vis_tbit_o));
assign Gwkiu6 = (Wxkiu6 & Dykiu6);
assign Dykiu6 = (Lm8iu6 | Kykiu6);
assign Wxkiu6 = (Hx9iu6 | Rykiu6);
assign Eashu6 = (Ydkiu6 ? Zvkiu6 : vis_psp_o[22]);
assign X9shu6 = (Fekiu6 ? Zvkiu6 : vis_msp_o[22]);
assign Q9shu6 = (Mekiu6 ? vis_r14_o[24] : Zvkiu6);
assign J9shu6 = (Tekiu6 ? vis_r12_o[24] : Zvkiu6);
assign C9shu6 = (Rdkiu6 ? vis_r7_o[24] : Zvkiu6);
assign V8shu6 = (Kdkiu6 ? vis_r6_o[24] : Zvkiu6);
assign O8shu6 = (Ddkiu6 ? vis_r5_o[24] : Zvkiu6);
assign H8shu6 = (Wckiu6 ? vis_r4_o[24] : Zvkiu6);
assign A8shu6 = (Afkiu6 ? vis_r11_o[24] : Zvkiu6);
assign T7shu6 = (Hfkiu6 ? vis_r10_o[24] : Zvkiu6);
assign M7shu6 = (Ofkiu6 ? vis_r9_o[24] : Zvkiu6);
assign F7shu6 = (Pckiu6 ? vis_r3_o[24] : Zvkiu6);
assign Y6shu6 = (Ickiu6 ? vis_r2_o[24] : Zvkiu6);
assign R6shu6 = (Mx8iu6 ? vis_r1_o[24] : Zvkiu6);
assign K6shu6 = (Lf8iu6 ? vis_r0_o[24] : Zvkiu6);
assign Zvkiu6 = (Nu8iu6 | Yykiu6);
assign D6shu6 = (Vfkiu6 ? vis_r8_o[26] : Fzkiu6);
assign W5shu6 = (~(Mzkiu6 & Tzkiu6));
assign Tzkiu6 = (A0liu6 & H0liu6);
assign H0liu6 = (~(Jl8iu6 & H0epw6));
assign A0liu6 = (~(vis_pc_o[25] & Ok8iu6));
assign Mzkiu6 = (O0liu6 & V0liu6);
assign V0liu6 = (~(W29iu6 & Fkfpw6[26]));
assign O0liu6 = (Hx9iu6 | C1liu6);
assign P5shu6 = (Ydkiu6 ? Fzkiu6 : vis_psp_o[24]);
assign I5shu6 = (Fekiu6 ? Fzkiu6 : vis_msp_o[24]);
assign B5shu6 = (Mekiu6 ? vis_r14_o[26] : Fzkiu6);
assign U4shu6 = (Tekiu6 ? vis_r12_o[26] : Fzkiu6);
assign N4shu6 = (Rdkiu6 ? vis_r7_o[26] : Fzkiu6);
assign G4shu6 = (Kdkiu6 ? vis_r6_o[26] : Fzkiu6);
assign Z3shu6 = (Ddkiu6 ? vis_r5_o[26] : Fzkiu6);
assign S3shu6 = (Wckiu6 ? vis_r4_o[26] : Fzkiu6);
assign L3shu6 = (Afkiu6 ? vis_r11_o[26] : Fzkiu6);
assign E3shu6 = (Hfkiu6 ? vis_r10_o[26] : Fzkiu6);
assign X2shu6 = (Ofkiu6 ? vis_r9_o[26] : Fzkiu6);
assign Q2shu6 = (Pckiu6 ? vis_r3_o[26] : Fzkiu6);
assign J2shu6 = (Ickiu6 ? vis_r2_o[26] : Fzkiu6);
assign C2shu6 = (Mx8iu6 ? vis_r1_o[26] : Fzkiu6);
assign V1shu6 = (Lf8iu6 ? vis_r0_o[26] : Fzkiu6);
assign Fzkiu6 = (J1liu6 | Q1liu6);
assign O1shu6 = (Vfkiu6 ? vis_r8_o[27] : X1liu6);
assign H1shu6 = (~(E2liu6 & L2liu6));
assign L2liu6 = (S2liu6 & Z2liu6);
assign Z2liu6 = (~(Jl8iu6 & O0epw6));
assign S2liu6 = (~(vis_pc_o[26] & Ok8iu6));
assign E2liu6 = (G3liu6 & N3liu6);
assign N3liu6 = (~(W29iu6 & Fkfpw6[27]));
assign G3liu6 = (Hx9iu6 | U3liu6);
assign A1shu6 = (Ydkiu6 ? X1liu6 : vis_psp_o[25]);
assign T0shu6 = (Fekiu6 ? X1liu6 : vis_msp_o[25]);
assign M0shu6 = (Mekiu6 ? vis_r14_o[27] : X1liu6);
assign F0shu6 = (Tekiu6 ? vis_r12_o[27] : X1liu6);
assign Yzrhu6 = (Rdkiu6 ? vis_r7_o[27] : X1liu6);
assign Rzrhu6 = (Kdkiu6 ? vis_r6_o[27] : X1liu6);
assign Kzrhu6 = (Ddkiu6 ? vis_r5_o[27] : X1liu6);
assign Dzrhu6 = (Wckiu6 ? vis_r4_o[27] : X1liu6);
assign Wyrhu6 = (Afkiu6 ? vis_r11_o[27] : X1liu6);
assign Pyrhu6 = (Hfkiu6 ? vis_r10_o[27] : X1liu6);
assign Iyrhu6 = (Ofkiu6 ? vis_r9_o[27] : X1liu6);
assign Byrhu6 = (Pckiu6 ? vis_r3_o[27] : X1liu6);
assign Uxrhu6 = (Ickiu6 ? vis_r2_o[27] : X1liu6);
assign Nxrhu6 = (Mx8iu6 ? vis_r1_o[27] : X1liu6);
assign Gxrhu6 = (Lf8iu6 ? vis_r0_o[27] : X1liu6);
assign X1liu6 = (B4liu6 | I4liu6);
assign Zwrhu6 = (Vfkiu6 ? vis_r8_o[29] : P4liu6);
assign Swrhu6 = (Ydkiu6 ? P4liu6 : vis_psp_o[27]);
assign Lwrhu6 = (Fekiu6 ? P4liu6 : vis_msp_o[27]);
assign Ewrhu6 = (Mekiu6 ? vis_r14_o[29] : P4liu6);
assign Xvrhu6 = (Tekiu6 ? vis_r12_o[29] : P4liu6);
assign Qvrhu6 = (Rdkiu6 ? vis_r7_o[29] : P4liu6);
assign Jvrhu6 = (Kdkiu6 ? vis_r6_o[29] : P4liu6);
assign Cvrhu6 = (Ddkiu6 ? vis_r5_o[29] : P4liu6);
assign Vurhu6 = (Wckiu6 ? vis_r4_o[29] : P4liu6);
assign Ourhu6 = (Afkiu6 ? vis_r11_o[29] : P4liu6);
assign Hurhu6 = (Hfkiu6 ? vis_r10_o[29] : P4liu6);
assign Aurhu6 = (Ofkiu6 ? vis_r9_o[29] : P4liu6);
assign Ttrhu6 = (Pckiu6 ? vis_r3_o[29] : P4liu6);
assign Mtrhu6 = (Ickiu6 ? vis_r2_o[29] : P4liu6);
assign Ftrhu6 = (Mx8iu6 ? vis_r1_o[29] : P4liu6);
assign Ysrhu6 = (Lf8iu6 ? vis_r0_o[29] : P4liu6);
assign P4liu6 = (Fj8iu6 | W4liu6);
assign Rsrhu6 = (Vfkiu6 ? vis_r8_o[30] : K39iu6);
assign K39iu6 = (~(D5liu6 & K5liu6));
assign Ksrhu6 = (Y5liu6 ? R5liu6 : vis_apsr_o[2]);
assign R5liu6 = (~(F6liu6 & M6liu6));
assign M6liu6 = (~(Ph8iu6 & T6liu6));
assign F6liu6 = (A7liu6 & H7liu6);
assign H7liu6 = (O7liu6 | V7liu6);
assign A7liu6 = (Cs8iu6 | D5liu6);
assign Dsrhu6 = (~(C8liu6 & J8liu6));
assign J8liu6 = (Q8liu6 & X8liu6);
assign X8liu6 = (~(Ok8iu6 & vis_pc_o[29]));
assign Q8liu6 = (E9liu6 & L9liu6);
assign L9liu6 = (~(Jl8iu6 & Rx0iu6));
assign E9liu6 = (~(vis_apsr_o[2] & Ql8iu6));
assign C8liu6 = (S9liu6 & Z9liu6);
assign Z9liu6 = (Lm8iu6 | Galiu6);
assign S9liu6 = (Hx9iu6 | Naliu6);
assign Wrrhu6 = (Vfkiu6 ? vis_r8_o[31] : D39iu6);
assign D39iu6 = (~(Ualiu6 & Bbliu6));
assign Prrhu6 = (Vfkiu6 ? vis_r8_o[0] : Tx8iu6);
assign Tx8iu6 = (~(Zt8iu6 & Ibliu6));
assign Zt8iu6 = (Pbliu6 & Wbliu6);
assign Wbliu6 = (Dcliu6 & Kcliu6);
assign Kcliu6 = (Rcliu6 | Ycliu6);
assign Dcliu6 = (Fdliu6 & Mdliu6);
assign Fdliu6 = (~(Tdliu6 & Aeliu6));
assign Pbliu6 = (Heliu6 & Oeliu6);
assign Oeliu6 = (Veliu6 | Cfliu6);
assign Heliu6 = (~(Jfliu6 & Qfliu6));
assign Irrhu6 = (~(Xfliu6 & Egliu6));
assign Egliu6 = (Lgliu6 & Sgliu6);
assign Sgliu6 = (~(Ok8iu6 & vis_pc_o[0]));
assign Lgliu6 = (Zgliu6 & Ghliu6);
assign Ghliu6 = (~(Nhliu6 & Uhliu6));
assign Uhliu6 = (Biliu6 & Iiliu6);
assign Nhliu6 = (Jl8iu6 & Piliu6);
assign Piliu6 = (Wiliu6 | Oviiu6);
assign Zgliu6 = (~(Ql8iu6 & vis_ipsr_o[1]));
assign Xfliu6 = (Djliu6 & Kjliu6);
assign Kjliu6 = (Lm8iu6 | Rjliu6);
assign Djliu6 = (Hx9iu6 | A34iu6);
assign Brrhu6 = (Fkliu6 ? Yjliu6 : vis_control_o);
assign Fkliu6 = (HREADY & Mkliu6);
assign Mkliu6 = (~(Tkliu6 & Alliu6));
assign Alliu6 = (~(Hlliu6 & Olliu6));
assign Olliu6 = (~(Vlliu6 & Cmliu6));
assign Cmliu6 = (~(Jmliu6 & S8fpw6[2]));
assign Jmliu6 = (S8fpw6[4] & Qmliu6);
assign Tkliu6 = (~(Clfiu6 | Xmliu6));
assign Yjliu6 = (~(Enliu6 & Lnliu6));
assign Lnliu6 = (~(Snliu6 & Qmliu6));
assign Snliu6 = (Wofiu6 ? Goliu6 : Znliu6);
assign Enliu6 = (Quzhu6 | Noliu6);
assign Uqrhu6 = (Mekiu6 ? vis_r14_o[1] : Uoliu6);
assign Nqrhu6 = (Tekiu6 ? vis_r12_o[1] : Uoliu6);
assign Gqrhu6 = (Rdkiu6 ? vis_r7_o[1] : Uoliu6);
assign Zprhu6 = (Kdkiu6 ? vis_r6_o[1] : Uoliu6);
assign Sprhu6 = (Ddkiu6 ? vis_r5_o[1] : Uoliu6);
assign Lprhu6 = (Wckiu6 ? vis_r4_o[1] : Uoliu6);
assign Eprhu6 = (Afkiu6 ? vis_r11_o[1] : Uoliu6);
assign Xorhu6 = (Hfkiu6 ? vis_r10_o[1] : Uoliu6);
assign Qorhu6 = (Ofkiu6 ? vis_r9_o[1] : Uoliu6);
assign Jorhu6 = (Vfkiu6 ? vis_r8_o[1] : Uoliu6);
assign Corhu6 = (Pckiu6 ? vis_r3_o[1] : Uoliu6);
assign Vnrhu6 = (Ickiu6 ? vis_r2_o[1] : Uoliu6);
assign Onrhu6 = (Mx8iu6 ? vis_r1_o[1] : Uoliu6);
assign Hnrhu6 = (Lf8iu6 ? vis_r0_o[1] : Uoliu6);
assign Uoliu6 = (~(Njciu6 & Bpliu6));
assign Anrhu6 = (~(Ipliu6 & Ppliu6));
assign Ppliu6 = (Wpliu6 & Dqliu6);
assign Dqliu6 = (~(vis_pc_o[24] & Ok8iu6));
assign Wpliu6 = (Kqliu6 & Rqliu6);
assign Rqliu6 = (~(vis_control_o & B29iu6));
assign B29iu6 = (Yqliu6 & Frliu6);
assign Yqliu6 = (~(U19iu6 | W29iu6));
assign Kqliu6 = (~(Jl8iu6 & A0epw6));
assign Ipliu6 = (Mrliu6 & Trliu6);
assign Trliu6 = (~(W29iu6 & Fkfpw6[25]));
assign Mrliu6 = (Hx9iu6 | Asliu6);
assign Tmrhu6 = (Ydkiu6 ? Hsliu6 : vis_psp_o[23]);
assign Mmrhu6 = (Fekiu6 ? Hsliu6 : vis_msp_o[23]);
assign Fmrhu6 = (Mekiu6 ? vis_r14_o[25] : Hsliu6);
assign Ylrhu6 = (Tekiu6 ? vis_r12_o[25] : Hsliu6);
assign Rlrhu6 = (Rdkiu6 ? vis_r7_o[25] : Hsliu6);
assign Klrhu6 = (Kdkiu6 ? vis_r6_o[25] : Hsliu6);
assign Dlrhu6 = (Ddkiu6 ? vis_r5_o[25] : Hsliu6);
assign Wkrhu6 = (Wckiu6 ? vis_r4_o[25] : Hsliu6);
assign Pkrhu6 = (Afkiu6 ? vis_r11_o[25] : Hsliu6);
assign Ikrhu6 = (Hfkiu6 ? vis_r10_o[25] : Hsliu6);
assign Bkrhu6 = (Ofkiu6 ? vis_r9_o[25] : Hsliu6);
assign Ujrhu6 = (Vfkiu6 ? vis_r8_o[25] : Hsliu6);
assign Njrhu6 = (Pckiu6 ? vis_r3_o[25] : Hsliu6);
assign Gjrhu6 = (Ickiu6 ? vis_r2_o[25] : Hsliu6);
assign Zirhu6 = (Mx8iu6 ? vis_r1_o[25] : Hsliu6);
assign Sirhu6 = (Lf8iu6 ? vis_r0_o[25] : Hsliu6);
assign Hsliu6 = (Osliu6 | Vsliu6);
assign Lirhu6 = (Hy8iu6 ? Iiliu6 : Iwfpw6[1]);
assign Hy8iu6 = (~(Eh6iu6 | L18iu6));
assign Eirhu6 = (~(Ctliu6 & Jtliu6));
assign Jtliu6 = (Qtliu6 & Xtliu6);
assign Xtliu6 = (~(Jl8iu6 & Fzdpw6));
assign Qtliu6 = (~(vis_pc_o[21] & Ok8iu6));
assign Ctliu6 = (Euliu6 & Luliu6);
assign Luliu6 = (Lm8iu6 | Suliu6);
assign Euliu6 = (~(Zm8iu6 & P74iu6));
assign Xhrhu6 = (Ydkiu6 ? Zuliu6 : vis_psp_o[20]);
assign Qhrhu6 = (Fekiu6 ? Zuliu6 : vis_msp_o[20]);
assign Jhrhu6 = (Mekiu6 ? vis_r14_o[22] : Zuliu6);
assign Chrhu6 = (Tekiu6 ? vis_r12_o[22] : Zuliu6);
assign Vgrhu6 = (Rdkiu6 ? vis_r7_o[22] : Zuliu6);
assign Ogrhu6 = (Kdkiu6 ? vis_r6_o[22] : Zuliu6);
assign Hgrhu6 = (Ddkiu6 ? vis_r5_o[22] : Zuliu6);
assign Agrhu6 = (Wckiu6 ? vis_r4_o[22] : Zuliu6);
assign Tfrhu6 = (Afkiu6 ? vis_r11_o[22] : Zuliu6);
assign Mfrhu6 = (Hfkiu6 ? vis_r10_o[22] : Zuliu6);
assign Ffrhu6 = (Ofkiu6 ? vis_r9_o[22] : Zuliu6);
assign Yerhu6 = (Vfkiu6 ? vis_r8_o[22] : Zuliu6);
assign Rerhu6 = (Pckiu6 ? vis_r3_o[22] : Zuliu6);
assign Kerhu6 = (Ickiu6 ? vis_r2_o[22] : Zuliu6);
assign Derhu6 = (Mx8iu6 ? vis_r1_o[22] : Zuliu6);
assign Wdrhu6 = (Lf8iu6 ? vis_r0_o[22] : Zuliu6);
assign Zuliu6 = (~(Gvliu6 & Nvliu6));
assign Gvliu6 = (Uvliu6 & Svkiu6);
assign Pdrhu6 = (~(Bwliu6 & Iwliu6));
assign Iwliu6 = (Pwliu6 & Wwliu6);
assign Wwliu6 = (~(Jl8iu6 & Yydpw6));
assign Pwliu6 = (~(vis_pc_o[20] & Ok8iu6));
assign Bwliu6 = (Dxliu6 & Kxliu6);
assign Kxliu6 = (Lm8iu6 | Rxliu6);
assign Dxliu6 = (Hx9iu6 | Yxliu6);
assign Idrhu6 = (Ydkiu6 ? Fyliu6 : vis_psp_o[19]);
assign Bdrhu6 = (Fekiu6 ? Fyliu6 : vis_msp_o[19]);
assign Ucrhu6 = (Mekiu6 ? vis_r14_o[21] : Fyliu6);
assign Ncrhu6 = (Tekiu6 ? vis_r12_o[21] : Fyliu6);
assign Gcrhu6 = (Rdkiu6 ? vis_r7_o[21] : Fyliu6);
assign Zbrhu6 = (Kdkiu6 ? vis_r6_o[21] : Fyliu6);
assign Sbrhu6 = (Ddkiu6 ? vis_r5_o[21] : Fyliu6);
assign Lbrhu6 = (Wckiu6 ? vis_r4_o[21] : Fyliu6);
assign Ebrhu6 = (Afkiu6 ? vis_r11_o[21] : Fyliu6);
assign Xarhu6 = (Hfkiu6 ? vis_r10_o[21] : Fyliu6);
assign Qarhu6 = (Ofkiu6 ? vis_r9_o[21] : Fyliu6);
assign Jarhu6 = (Vfkiu6 ? vis_r8_o[21] : Fyliu6);
assign Carhu6 = (Pckiu6 ? vis_r3_o[21] : Fyliu6);
assign V9rhu6 = (Ickiu6 ? vis_r2_o[21] : Fyliu6);
assign O9rhu6 = (Mx8iu6 ? vis_r1_o[21] : Fyliu6);
assign H9rhu6 = (Lf8iu6 ? vis_r0_o[21] : Fyliu6);
assign Fyliu6 = (~(Myliu6 & Tyliu6));
assign Myliu6 = (Azliu6 & Svkiu6);
assign A9rhu6 = (~(Hzliu6 & Ozliu6));
assign Ozliu6 = (Vzliu6 & C0miu6);
assign C0miu6 = (~(Jl8iu6 & Rydpw6));
assign Vzliu6 = (~(vis_pc_o[19] & Ok8iu6));
assign Hzliu6 = (J0miu6 & Q0miu6);
assign Q0miu6 = (Lm8iu6 | X0miu6);
assign J0miu6 = (~(Zm8iu6 & B74iu6));
assign T8rhu6 = (Ydkiu6 ? E1miu6 : vis_psp_o[18]);
assign M8rhu6 = (Fekiu6 ? E1miu6 : vis_msp_o[18]);
assign F8rhu6 = (Mekiu6 ? vis_r14_o[20] : E1miu6);
assign Y7rhu6 = (Tekiu6 ? vis_r12_o[20] : E1miu6);
assign R7rhu6 = (Rdkiu6 ? vis_r7_o[20] : E1miu6);
assign K7rhu6 = (Kdkiu6 ? vis_r6_o[20] : E1miu6);
assign D7rhu6 = (Ddkiu6 ? vis_r5_o[20] : E1miu6);
assign W6rhu6 = (Wckiu6 ? vis_r4_o[20] : E1miu6);
assign P6rhu6 = (Afkiu6 ? vis_r11_o[20] : E1miu6);
assign I6rhu6 = (Hfkiu6 ? vis_r10_o[20] : E1miu6);
assign B6rhu6 = (Ofkiu6 ? vis_r9_o[20] : E1miu6);
assign U5rhu6 = (Vfkiu6 ? vis_r8_o[20] : E1miu6);
assign N5rhu6 = (Pckiu6 ? vis_r3_o[20] : E1miu6);
assign G5rhu6 = (Ickiu6 ? vis_r2_o[20] : E1miu6);
assign Z4rhu6 = (Mx8iu6 ? vis_r1_o[20] : E1miu6);
assign S4rhu6 = (Lf8iu6 ? vis_r0_o[20] : E1miu6);
assign E1miu6 = (~(L1miu6 & S1miu6));
assign L1miu6 = (Z1miu6 & Svkiu6);
assign L4rhu6 = (~(G2miu6 & N2miu6));
assign N2miu6 = (U2miu6 & B3miu6);
assign B3miu6 = (~(Jl8iu6 & Kydpw6));
assign U2miu6 = (~(vis_pc_o[18] & Ok8iu6));
assign G2miu6 = (I3miu6 & P3miu6);
assign P3miu6 = (Lm8iu6 | W3miu6);
assign I3miu6 = (~(Zm8iu6 & U64iu6));
assign E4rhu6 = (Ydkiu6 ? D4miu6 : vis_psp_o[17]);
assign X3rhu6 = (Fekiu6 ? D4miu6 : vis_msp_o[17]);
assign Q3rhu6 = (Mekiu6 ? vis_r14_o[19] : D4miu6);
assign J3rhu6 = (Tekiu6 ? vis_r12_o[19] : D4miu6);
assign C3rhu6 = (Rdkiu6 ? vis_r7_o[19] : D4miu6);
assign V2rhu6 = (Kdkiu6 ? vis_r6_o[19] : D4miu6);
assign O2rhu6 = (Ddkiu6 ? vis_r5_o[19] : D4miu6);
assign H2rhu6 = (Wckiu6 ? vis_r4_o[19] : D4miu6);
assign A2rhu6 = (Afkiu6 ? vis_r11_o[19] : D4miu6);
assign T1rhu6 = (Hfkiu6 ? vis_r10_o[19] : D4miu6);
assign M1rhu6 = (Ofkiu6 ? vis_r9_o[19] : D4miu6);
assign F1rhu6 = (Vfkiu6 ? vis_r8_o[19] : D4miu6);
assign Y0rhu6 = (Pckiu6 ? vis_r3_o[19] : D4miu6);
assign R0rhu6 = (Ickiu6 ? vis_r2_o[19] : D4miu6);
assign K0rhu6 = (Mx8iu6 ? vis_r1_o[19] : D4miu6);
assign D0rhu6 = (Lf8iu6 ? vis_r0_o[19] : D4miu6);
assign D4miu6 = (~(K4miu6 & R4miu6));
assign K4miu6 = (Y4miu6 & Svkiu6);
assign Wzqhu6 = (~(F5miu6 & M5miu6));
assign M5miu6 = (T5miu6 & A6miu6);
assign A6miu6 = (~(Jl8iu6 & Dydpw6));
assign T5miu6 = (~(vis_pc_o[17] & Ok8iu6));
assign F5miu6 = (H6miu6 & O6miu6);
assign O6miu6 = (Lm8iu6 | V6miu6);
assign H6miu6 = (~(Zm8iu6 & N64iu6));
assign Pzqhu6 = (Ydkiu6 ? C7miu6 : vis_psp_o[16]);
assign Izqhu6 = (Fekiu6 ? C7miu6 : vis_msp_o[16]);
assign Bzqhu6 = (Mekiu6 ? vis_r14_o[18] : C7miu6);
assign Uyqhu6 = (Tekiu6 ? vis_r12_o[18] : C7miu6);
assign Nyqhu6 = (Rdkiu6 ? vis_r7_o[18] : C7miu6);
assign Gyqhu6 = (Kdkiu6 ? vis_r6_o[18] : C7miu6);
assign Zxqhu6 = (Ddkiu6 ? vis_r5_o[18] : C7miu6);
assign Sxqhu6 = (Wckiu6 ? vis_r4_o[18] : C7miu6);
assign Lxqhu6 = (Afkiu6 ? vis_r11_o[18] : C7miu6);
assign Exqhu6 = (Hfkiu6 ? vis_r10_o[18] : C7miu6);
assign Xwqhu6 = (Ofkiu6 ? vis_r9_o[18] : C7miu6);
assign Qwqhu6 = (Vfkiu6 ? vis_r8_o[18] : C7miu6);
assign Jwqhu6 = (Pckiu6 ? vis_r3_o[18] : C7miu6);
assign Cwqhu6 = (Ickiu6 ? vis_r2_o[18] : C7miu6);
assign Vvqhu6 = (Mx8iu6 ? vis_r1_o[18] : C7miu6);
assign Ovqhu6 = (Lf8iu6 ? vis_r0_o[18] : C7miu6);
assign C7miu6 = (~(J7miu6 & Q7miu6));
assign J7miu6 = (X7miu6 & Svkiu6);
assign Hvqhu6 = (~(E8miu6 & L8miu6));
assign L8miu6 = (S8miu6 & Z8miu6);
assign Z8miu6 = (~(Jl8iu6 & Wxdpw6));
assign S8miu6 = (~(vis_pc_o[16] & Ok8iu6));
assign E8miu6 = (G9miu6 & N9miu6);
assign N9miu6 = (Lm8iu6 | U9miu6);
assign G9miu6 = (~(Zm8iu6 & G64iu6));
assign Avqhu6 = (Ydkiu6 ? Bamiu6 : vis_psp_o[15]);
assign Tuqhu6 = (Fekiu6 ? Bamiu6 : vis_msp_o[15]);
assign Muqhu6 = (Mekiu6 ? vis_r14_o[17] : Bamiu6);
assign Fuqhu6 = (Tekiu6 ? vis_r12_o[17] : Bamiu6);
assign Ytqhu6 = (Rdkiu6 ? vis_r7_o[17] : Bamiu6);
assign Rtqhu6 = (Kdkiu6 ? vis_r6_o[17] : Bamiu6);
assign Ktqhu6 = (Ddkiu6 ? vis_r5_o[17] : Bamiu6);
assign Dtqhu6 = (Wckiu6 ? vis_r4_o[17] : Bamiu6);
assign Wsqhu6 = (Afkiu6 ? vis_r11_o[17] : Bamiu6);
assign Psqhu6 = (Hfkiu6 ? vis_r10_o[17] : Bamiu6);
assign Isqhu6 = (Ofkiu6 ? vis_r9_o[17] : Bamiu6);
assign Bsqhu6 = (Vfkiu6 ? vis_r8_o[17] : Bamiu6);
assign Urqhu6 = (Pckiu6 ? vis_r3_o[17] : Bamiu6);
assign Nrqhu6 = (Ickiu6 ? vis_r2_o[17] : Bamiu6);
assign Grqhu6 = (Mx8iu6 ? vis_r1_o[17] : Bamiu6);
assign Zqqhu6 = (Lf8iu6 ? vis_r0_o[17] : Bamiu6);
assign Bamiu6 = (~(Iamiu6 & Pamiu6));
assign Iamiu6 = (Wamiu6 & Svkiu6);
assign Sqqhu6 = (~(Dbmiu6 & Kbmiu6));
assign Kbmiu6 = (Rbmiu6 & Ybmiu6);
assign Ybmiu6 = (~(Jl8iu6 & Pxdpw6));
assign Rbmiu6 = (~(vis_pc_o[15] & Ok8iu6));
assign Dbmiu6 = (Fcmiu6 & Mcmiu6);
assign Mcmiu6 = (Lm8iu6 | Tcmiu6);
assign Fcmiu6 = (~(Zm8iu6 & Z54iu6));
assign Lqqhu6 = (Ydkiu6 ? Admiu6 : vis_psp_o[14]);
assign Eqqhu6 = (Fekiu6 ? Admiu6 : vis_msp_o[14]);
assign Xpqhu6 = (Mekiu6 ? vis_r14_o[16] : Admiu6);
assign Qpqhu6 = (Tekiu6 ? vis_r12_o[16] : Admiu6);
assign Jpqhu6 = (Rdkiu6 ? vis_r7_o[16] : Admiu6);
assign Cpqhu6 = (Kdkiu6 ? vis_r6_o[16] : Admiu6);
assign Voqhu6 = (Ddkiu6 ? vis_r5_o[16] : Admiu6);
assign Ooqhu6 = (Wckiu6 ? vis_r4_o[16] : Admiu6);
assign Hoqhu6 = (Afkiu6 ? vis_r11_o[16] : Admiu6);
assign Aoqhu6 = (Hfkiu6 ? vis_r10_o[16] : Admiu6);
assign Tnqhu6 = (Ofkiu6 ? vis_r9_o[16] : Admiu6);
assign Mnqhu6 = (Vfkiu6 ? vis_r8_o[16] : Admiu6);
assign Fnqhu6 = (Pckiu6 ? vis_r3_o[16] : Admiu6);
assign Ymqhu6 = (Ickiu6 ? vis_r2_o[16] : Admiu6);
assign Rmqhu6 = (Mx8iu6 ? vis_r1_o[16] : Admiu6);
assign Kmqhu6 = (Lf8iu6 ? vis_r0_o[16] : Admiu6);
assign Admiu6 = (~(Hdmiu6 & Odmiu6));
assign Hdmiu6 = (Vdmiu6 & Svkiu6);
assign Dmqhu6 = (~(Cemiu6 & Jemiu6));
assign Jemiu6 = (Qemiu6 & Xemiu6);
assign Xemiu6 = (~(Jl8iu6 & Tugpw6[13]));
assign Qemiu6 = (~(vis_pc_o[14] & Ok8iu6));
assign Cemiu6 = (Efmiu6 & Lfmiu6);
assign Lfmiu6 = (Lm8iu6 | Sfmiu6);
assign Efmiu6 = (~(Zm8iu6 & S54iu6));
assign Wlqhu6 = (Ydkiu6 ? Zfmiu6 : vis_psp_o[13]);
assign Plqhu6 = (Fekiu6 ? Zfmiu6 : vis_msp_o[13]);
assign Ilqhu6 = (Mekiu6 ? vis_r14_o[15] : Zfmiu6);
assign Blqhu6 = (Tekiu6 ? vis_r12_o[15] : Zfmiu6);
assign Ukqhu6 = (Rdkiu6 ? vis_r7_o[15] : Zfmiu6);
assign Nkqhu6 = (Kdkiu6 ? vis_r6_o[15] : Zfmiu6);
assign Gkqhu6 = (Ddkiu6 ? vis_r5_o[15] : Zfmiu6);
assign Zjqhu6 = (Wckiu6 ? vis_r4_o[15] : Zfmiu6);
assign Sjqhu6 = (Afkiu6 ? vis_r11_o[15] : Zfmiu6);
assign Ljqhu6 = (Hfkiu6 ? vis_r10_o[15] : Zfmiu6);
assign Ejqhu6 = (Ofkiu6 ? vis_r9_o[15] : Zfmiu6);
assign Xiqhu6 = (Vfkiu6 ? vis_r8_o[15] : Zfmiu6);
assign Qiqhu6 = (Pckiu6 ? vis_r3_o[15] : Zfmiu6);
assign Jiqhu6 = (Ickiu6 ? vis_r2_o[15] : Zfmiu6);
assign Ciqhu6 = (Mx8iu6 ? vis_r1_o[15] : Zfmiu6);
assign Vhqhu6 = (Lf8iu6 ? vis_r0_o[15] : Zfmiu6);
assign Zfmiu6 = (~(Ggmiu6 & Ngmiu6));
assign Ohqhu6 = (~(Ugmiu6 & Bhmiu6));
assign Bhmiu6 = (Ihmiu6 & Phmiu6);
assign Phmiu6 = (~(Jl8iu6 & Tugpw6[12]));
assign Ihmiu6 = (~(vis_pc_o[13] & Ok8iu6));
assign Ugmiu6 = (Whmiu6 & Dimiu6);
assign Dimiu6 = (Lm8iu6 | Kimiu6);
assign Whmiu6 = (~(Zm8iu6 & L54iu6));
assign Hhqhu6 = (Ydkiu6 ? Rimiu6 : vis_psp_o[12]);
assign Ahqhu6 = (Fekiu6 ? Rimiu6 : vis_msp_o[12]);
assign Tgqhu6 = (Mekiu6 ? vis_r14_o[14] : Rimiu6);
assign Mgqhu6 = (Tekiu6 ? vis_r12_o[14] : Rimiu6);
assign Fgqhu6 = (Rdkiu6 ? vis_r7_o[14] : Rimiu6);
assign Yfqhu6 = (Kdkiu6 ? vis_r6_o[14] : Rimiu6);
assign Rfqhu6 = (Ddkiu6 ? vis_r5_o[14] : Rimiu6);
assign Kfqhu6 = (Wckiu6 ? vis_r4_o[14] : Rimiu6);
assign Dfqhu6 = (Afkiu6 ? vis_r11_o[14] : Rimiu6);
assign Weqhu6 = (Hfkiu6 ? vis_r10_o[14] : Rimiu6);
assign Peqhu6 = (Ofkiu6 ? vis_r9_o[14] : Rimiu6);
assign Ieqhu6 = (Vfkiu6 ? vis_r8_o[14] : Rimiu6);
assign Beqhu6 = (Pckiu6 ? vis_r3_o[14] : Rimiu6);
assign Udqhu6 = (Ickiu6 ? vis_r2_o[14] : Rimiu6);
assign Ndqhu6 = (Mx8iu6 ? vis_r1_o[14] : Rimiu6);
assign Gdqhu6 = (Lf8iu6 ? vis_r0_o[14] : Rimiu6);
assign Rimiu6 = (Yimiu6 | Fjmiu6);
assign Zcqhu6 = (~(Mjmiu6 & Tjmiu6));
assign Tjmiu6 = (Akmiu6 & Hkmiu6);
assign Hkmiu6 = (~(Jl8iu6 & Tugpw6[11]));
assign Akmiu6 = (~(vis_pc_o[12] & Ok8iu6));
assign Mjmiu6 = (Okmiu6 & Vkmiu6);
assign Vkmiu6 = (Lm8iu6 | Clmiu6);
assign Okmiu6 = (~(Zm8iu6 & E54iu6));
assign Scqhu6 = (Ydkiu6 ? Jlmiu6 : vis_psp_o[11]);
assign Lcqhu6 = (Fekiu6 ? Jlmiu6 : vis_msp_o[11]);
assign Ecqhu6 = (Mekiu6 ? vis_r14_o[13] : Jlmiu6);
assign Xbqhu6 = (Tekiu6 ? vis_r12_o[13] : Jlmiu6);
assign Qbqhu6 = (Rdkiu6 ? vis_r7_o[13] : Jlmiu6);
assign Jbqhu6 = (Kdkiu6 ? vis_r6_o[13] : Jlmiu6);
assign Cbqhu6 = (Ddkiu6 ? vis_r5_o[13] : Jlmiu6);
assign Vaqhu6 = (Wckiu6 ? vis_r4_o[13] : Jlmiu6);
assign Oaqhu6 = (Afkiu6 ? vis_r11_o[13] : Jlmiu6);
assign Haqhu6 = (Hfkiu6 ? vis_r10_o[13] : Jlmiu6);
assign Aaqhu6 = (Ofkiu6 ? vis_r9_o[13] : Jlmiu6);
assign T9qhu6 = (Vfkiu6 ? vis_r8_o[13] : Jlmiu6);
assign M9qhu6 = (Pckiu6 ? vis_r3_o[13] : Jlmiu6);
assign F9qhu6 = (Ickiu6 ? vis_r2_o[13] : Jlmiu6);
assign Y8qhu6 = (Mx8iu6 ? vis_r1_o[13] : Jlmiu6);
assign R8qhu6 = (Lf8iu6 ? vis_r0_o[13] : Jlmiu6);
assign Jlmiu6 = (Qlmiu6 | Xlmiu6);
assign K8qhu6 = (~(Emmiu6 & Lmmiu6));
assign Lmmiu6 = (Smmiu6 & Zmmiu6);
assign Zmmiu6 = (~(Jl8iu6 & Ixdpw6));
assign Smmiu6 = (~(vis_pc_o[11] & Ok8iu6));
assign Emmiu6 = (Gnmiu6 & Nnmiu6);
assign Nnmiu6 = (Lm8iu6 | Unmiu6);
assign Gnmiu6 = (~(Zm8iu6 & X44iu6));
assign D8qhu6 = (Ydkiu6 ? Bomiu6 : vis_psp_o[10]);
assign W7qhu6 = (Fekiu6 ? Bomiu6 : vis_msp_o[10]);
assign P7qhu6 = (Mekiu6 ? vis_r14_o[12] : Bomiu6);
assign I7qhu6 = (Tekiu6 ? vis_r12_o[12] : Bomiu6);
assign B7qhu6 = (Rdkiu6 ? vis_r7_o[12] : Bomiu6);
assign U6qhu6 = (Kdkiu6 ? vis_r6_o[12] : Bomiu6);
assign N6qhu6 = (Ddkiu6 ? vis_r5_o[12] : Bomiu6);
assign G6qhu6 = (Wckiu6 ? vis_r4_o[12] : Bomiu6);
assign Z5qhu6 = (Afkiu6 ? vis_r11_o[12] : Bomiu6);
assign S5qhu6 = (Hfkiu6 ? vis_r10_o[12] : Bomiu6);
assign L5qhu6 = (Ofkiu6 ? vis_r9_o[12] : Bomiu6);
assign E5qhu6 = (Vfkiu6 ? vis_r8_o[12] : Bomiu6);
assign X4qhu6 = (Pckiu6 ? vis_r3_o[12] : Bomiu6);
assign Q4qhu6 = (Ickiu6 ? vis_r2_o[12] : Bomiu6);
assign J4qhu6 = (Mx8iu6 ? vis_r1_o[12] : Bomiu6);
assign C4qhu6 = (Lf8iu6 ? vis_r0_o[12] : Bomiu6);
assign Bomiu6 = (Iomiu6 | Pomiu6);
assign V3qhu6 = (~(Womiu6 & Dpmiu6));
assign Dpmiu6 = (Kpmiu6 & Rpmiu6);
assign Rpmiu6 = (~(Jl8iu6 & Tugpw6[9]));
assign Tugpw6[9] = (~(Ypmiu6 & Fqmiu6));
assign Fqmiu6 = (~(N5fpw6[10] & Sdaiu6));
assign Ypmiu6 = (Mqmiu6 & Tqmiu6);
assign Tqmiu6 = (T2iiu6 | Sn0iu6);
assign Mqmiu6 = (~(Eafpw6[11] & A3iiu6));
assign Kpmiu6 = (~(vis_pc_o[10] & Ok8iu6));
assign Womiu6 = (Armiu6 & Hrmiu6);
assign Hrmiu6 = (Lm8iu6 | Ormiu6);
assign Armiu6 = (~(Zm8iu6 & Q44iu6));
assign O3qhu6 = (Ydkiu6 ? Vrmiu6 : vis_psp_o[9]);
assign H3qhu6 = (Fekiu6 ? Vrmiu6 : vis_msp_o[9]);
assign A3qhu6 = (Mekiu6 ? vis_r14_o[11] : Vrmiu6);
assign T2qhu6 = (Tekiu6 ? vis_r12_o[11] : Vrmiu6);
assign Tekiu6 = (!Csmiu6);
assign M2qhu6 = (Rdkiu6 ? vis_r7_o[11] : Vrmiu6);
assign Rdkiu6 = (!Jsmiu6);
assign F2qhu6 = (Kdkiu6 ? vis_r6_o[11] : Vrmiu6);
assign Y1qhu6 = (Ddkiu6 ? vis_r5_o[11] : Vrmiu6);
assign Ddkiu6 = (!Qsmiu6);
assign R1qhu6 = (Wckiu6 ? vis_r4_o[11] : Vrmiu6);
assign Wckiu6 = (!Xsmiu6);
assign K1qhu6 = (Afkiu6 ? vis_r11_o[11] : Vrmiu6);
assign Afkiu6 = (!Etmiu6);
assign D1qhu6 = (Hfkiu6 ? vis_r10_o[11] : Vrmiu6);
assign W0qhu6 = (Ofkiu6 ? vis_r9_o[11] : Vrmiu6);
assign Ofkiu6 = (!Ltmiu6);
assign P0qhu6 = (Vfkiu6 ? vis_r8_o[11] : Vrmiu6);
assign Vfkiu6 = (!Stmiu6);
assign I0qhu6 = (Pckiu6 ? vis_r3_o[11] : Vrmiu6);
assign Pckiu6 = (!Ztmiu6);
assign B0qhu6 = (Ickiu6 ? vis_r2_o[11] : Vrmiu6);
assign Uzphu6 = (Mx8iu6 ? vis_r1_o[11] : Vrmiu6);
assign Mx8iu6 = (!Gumiu6);
assign Nzphu6 = (Lf8iu6 ? vis_r0_o[11] : Vrmiu6);
assign Lf8iu6 = (!Numiu6);
assign Vrmiu6 = (Uumiu6 | Bvmiu6);
assign Gzphu6 = (~(Ivmiu6 & Pvmiu6));
assign Pvmiu6 = (Wvmiu6 & Dwmiu6);
assign Dwmiu6 = (~(Jl8iu6 & Tugpw6[8]));
assign Tugpw6[8] = (~(Kwmiu6 & Rwmiu6));
assign Rwmiu6 = (~(N5fpw6[9] & Sdaiu6));
assign Kwmiu6 = (Ywmiu6 & Fxmiu6);
assign Fxmiu6 = (T2iiu6 | Zn0iu6);
assign Ywmiu6 = (~(Eafpw6[10] & A3iiu6));
assign Wvmiu6 = (~(vis_pc_o[9] & Ok8iu6));
assign Ivmiu6 = (Mxmiu6 & Txmiu6);
assign Txmiu6 = (Lm8iu6 | Aymiu6);
assign Mxmiu6 = (~(Zm8iu6 & J44iu6));
assign Zyphu6 = (Ydkiu6 ? Hymiu6 : vis_psp_o[8]);
assign Syphu6 = (Fekiu6 ? Hymiu6 : vis_msp_o[8]);
assign Lyphu6 = (Mekiu6 ? vis_r14_o[10] : Hymiu6);
assign Eyphu6 = (Csmiu6 ? Hymiu6 : vis_r12_o[10]);
assign Xxphu6 = (Jsmiu6 ? Hymiu6 : vis_r7_o[10]);
assign Qxphu6 = (Kdkiu6 ? vis_r6_o[10] : Hymiu6);
assign Jxphu6 = (Qsmiu6 ? Hymiu6 : vis_r5_o[10]);
assign Cxphu6 = (Xsmiu6 ? Hymiu6 : vis_r4_o[10]);
assign Vwphu6 = (Etmiu6 ? Hymiu6 : vis_r11_o[10]);
assign Owphu6 = (Hfkiu6 ? vis_r10_o[10] : Hymiu6);
assign Hwphu6 = (Ltmiu6 ? Hymiu6 : vis_r9_o[10]);
assign Awphu6 = (Stmiu6 ? Hymiu6 : vis_r8_o[10]);
assign Tvphu6 = (Ztmiu6 ? Hymiu6 : vis_r3_o[10]);
assign Mvphu6 = (Ickiu6 ? vis_r2_o[10] : Hymiu6);
assign Fvphu6 = (Gumiu6 ? Hymiu6 : vis_r1_o[10]);
assign Yuphu6 = (Numiu6 ? Hymiu6 : vis_r0_o[10]);
assign Hymiu6 = (Oymiu6 | Vymiu6);
assign Ruphu6 = (Jzmiu6 ? Czmiu6 : L8ehu6);
assign Jzmiu6 = (Qzmiu6 & HREADY);
assign Qzmiu6 = (Xzmiu6 & E0niu6);
assign E0niu6 = (L0niu6 | Bi0iu6);
assign Czmiu6 = (Uzaiu6 ? Gh0iu6 : S0niu6);
assign Kuphu6 = (~(Z0niu6 & G1niu6));
assign G1niu6 = (N1niu6 & U1niu6);
assign U1niu6 = (~(vis_pc_o[8] & Ok8iu6));
assign N1niu6 = (B2niu6 & I2niu6);
assign I2niu6 = (~(P2niu6 & L8ehu6));
assign P2niu6 = (Ql8iu6 & Gc5iu6);
assign B2niu6 = (~(Jl8iu6 & Tugpw6[7]));
assign Z0niu6 = (W2niu6 & D3niu6);
assign D3niu6 = (~(W29iu6 & Fkfpw6[9]));
assign W2niu6 = (~(Zm8iu6 & Ym4iu6));
assign Duphu6 = (Ydkiu6 ? K3niu6 : vis_psp_o[7]);
assign Wtphu6 = (Fekiu6 ? K3niu6 : vis_msp_o[7]);
assign Ptphu6 = (Mekiu6 ? vis_r14_o[9] : K3niu6);
assign Itphu6 = (Csmiu6 ? K3niu6 : vis_r12_o[9]);
assign Btphu6 = (Jsmiu6 ? K3niu6 : vis_r7_o[9]);
assign Usphu6 = (Kdkiu6 ? vis_r6_o[9] : K3niu6);
assign Nsphu6 = (Qsmiu6 ? K3niu6 : vis_r5_o[9]);
assign Gsphu6 = (Xsmiu6 ? K3niu6 : vis_r4_o[9]);
assign Zrphu6 = (Etmiu6 ? K3niu6 : vis_r11_o[9]);
assign Srphu6 = (Hfkiu6 ? vis_r10_o[9] : K3niu6);
assign Lrphu6 = (Ltmiu6 ? K3niu6 : vis_r9_o[9]);
assign Erphu6 = (Stmiu6 ? K3niu6 : vis_r8_o[9]);
assign Xqphu6 = (Ztmiu6 ? K3niu6 : vis_r3_o[9]);
assign Qqphu6 = (Ickiu6 ? vis_r2_o[9] : K3niu6);
assign Jqphu6 = (Gumiu6 ? K3niu6 : vis_r1_o[9]);
assign Cqphu6 = (Numiu6 ? K3niu6 : vis_r0_o[9]);
assign K3niu6 = (S0niu6 | R3niu6);
assign Vpphu6 = (~(Y3niu6 & F4niu6));
assign F4niu6 = (M4niu6 & T4niu6);
assign T4niu6 = (~(Jl8iu6 & Tugpw6[6]));
assign Tugpw6[6] = (~(A5niu6 & H5niu6));
assign H5niu6 = (~(N5fpw6[7] & Sdaiu6));
assign A5niu6 = (O5niu6 & V5niu6);
assign V5niu6 = (T2iiu6 | Ve0iu6);
assign O5niu6 = (~(Eafpw6[8] & A3iiu6));
assign M4niu6 = (~(vis_pc_o[7] & Ok8iu6));
assign Y3niu6 = (C6niu6 & J6niu6);
assign J6niu6 = (Lm8iu6 | Q6niu6);
assign C6niu6 = (~(Zm8iu6 & Pl4iu6));
assign Opphu6 = (Ydkiu6 ? X6niu6 : vis_psp_o[6]);
assign Hpphu6 = (Fekiu6 ? X6niu6 : vis_msp_o[6]);
assign Apphu6 = (Mekiu6 ? vis_r14_o[8] : X6niu6);
assign Tophu6 = (Csmiu6 ? X6niu6 : vis_r12_o[8]);
assign Mophu6 = (Jsmiu6 ? X6niu6 : vis_r7_o[8]);
assign Fophu6 = (Kdkiu6 ? vis_r6_o[8] : X6niu6);
assign Ynphu6 = (Qsmiu6 ? X6niu6 : vis_r5_o[8]);
assign Rnphu6 = (Xsmiu6 ? X6niu6 : vis_r4_o[8]);
assign Knphu6 = (Etmiu6 ? X6niu6 : vis_r11_o[8]);
assign Dnphu6 = (Hfkiu6 ? vis_r10_o[8] : X6niu6);
assign Wmphu6 = (Ltmiu6 ? X6niu6 : vis_r9_o[8]);
assign Pmphu6 = (Stmiu6 ? X6niu6 : vis_r8_o[8]);
assign Imphu6 = (Ztmiu6 ? X6niu6 : vis_r3_o[8]);
assign Bmphu6 = (Ickiu6 ? vis_r2_o[8] : X6niu6);
assign Ulphu6 = (Gumiu6 ? X6niu6 : vis_r1_o[8]);
assign Nlphu6 = (Numiu6 ? X6niu6 : vis_r0_o[8]);
assign X6niu6 = (E7niu6 | L7niu6);
assign Glphu6 = (~(S7niu6 & Z7niu6));
assign Z7niu6 = (~(G8niu6 & Ug8iu6));
assign S7niu6 = (HREADY ? U8niu6 : N8niu6);
assign U8niu6 = (~(B9niu6 & I9niu6));
assign I9niu6 = (~(P9niu6 & Ug8iu6));
assign B9niu6 = (Ug8iu6 ? Daniu6 : W9niu6);
assign Daniu6 = (Kaniu6 & Raniu6);
assign Raniu6 = (~(Idfpw6[31] & Eafpw6[31]));
assign Kaniu6 = (D5epw6 ? Idfpw6[31] : Eafpw6[31]);
assign W9niu6 = (Yaniu6 & Fbniu6);
assign Fbniu6 = (~(Mbniu6 & Tbniu6));
assign Tbniu6 = (Cs8iu6 | Acniu6);
assign Yaniu6 = (~(Acniu6 & Hcniu6));
assign N8niu6 = (!vis_apsr_o[0]);
assign Zkphu6 = (~(Ocniu6 & Vcniu6));
assign Vcniu6 = (Cdniu6 & Jdniu6);
assign Jdniu6 = (~(Ok8iu6 & vis_pc_o[27]));
assign Cdniu6 = (Qdniu6 & Xdniu6);
assign Xdniu6 = (~(Jl8iu6 & V0epw6));
assign Qdniu6 = (~(vis_apsr_o[0] & Ql8iu6));
assign Ocniu6 = (Eeniu6 & Leniu6);
assign Leniu6 = (Lm8iu6 | Seniu6);
assign Eeniu6 = (Hx9iu6 | Zeniu6);
assign Skphu6 = (Ydkiu6 ? Gfniu6 : vis_psp_o[26]);
assign Ydkiu6 = (Nfniu6 & Vrfhu6);
assign Nfniu6 = (!Ufniu6);
assign Lkphu6 = (Fekiu6 ? Gfniu6 : vis_msp_o[26]);
assign Fekiu6 = (~(Ufniu6 | Vrfhu6));
assign Ufniu6 = (~(Bgniu6 & Igniu6));
assign Bgniu6 = (~(Pgniu6 | Wgniu6));
assign Ekphu6 = (Mekiu6 ? vis_r14_o[28] : Gfniu6);
assign Mekiu6 = (~(Dhniu6 & Khniu6));
assign Xjphu6 = (Csmiu6 ? Gfniu6 : vis_r12_o[28]);
assign Csmiu6 = (Rhniu6 & Khniu6);
assign Rhniu6 = (~(Yhniu6 | Wgniu6));
assign Qjphu6 = (Jsmiu6 ? Gfniu6 : vis_r7_o[28]);
assign Jsmiu6 = (Finiu6 & Miniu6);
assign Finiu6 = (Tiniu6 & Ajniu6);
assign Jjphu6 = (Kdkiu6 ? vis_r6_o[28] : Gfniu6);
assign Kdkiu6 = (~(Khniu6 & Miniu6));
assign Cjphu6 = (Qsmiu6 ? Gfniu6 : vis_r5_o[28]);
assign Qsmiu6 = (Hjniu6 & Igniu6);
assign Hjniu6 = (~(Ojniu6 | Pgniu6));
assign Viphu6 = (Xsmiu6 ? Gfniu6 : vis_r4_o[28]);
assign Xsmiu6 = (Vjniu6 & Khniu6);
assign Khniu6 = (~(Ajniu6 | Pgniu6));
assign Vjniu6 = (~(Yhniu6 | Ojniu6));
assign Oiphu6 = (Etmiu6 ? Gfniu6 : vis_r11_o[28]);
assign Etmiu6 = (Ckniu6 & Dhniu6);
assign Hiphu6 = (Hfkiu6 ? vis_r10_o[28] : Gfniu6);
assign Hfkiu6 = (~(Dhniu6 & Jkniu6));
assign Dhniu6 = (~(Wgniu6 | Qkniu6));
assign Aiphu6 = (Ltmiu6 ? Gfniu6 : vis_r9_o[28]);
assign Ltmiu6 = (Xkniu6 & Igniu6);
assign Xkniu6 = (~(Tiniu6 | Wgniu6));
assign Thphu6 = (Stmiu6 ? Gfniu6 : vis_r8_o[28]);
assign Stmiu6 = (Elniu6 & Qkniu6);
assign Elniu6 = (Jkniu6 & Ojniu6);
assign Mhphu6 = (Ztmiu6 ? Gfniu6 : vis_r3_o[28]);
assign Ztmiu6 = (Ckniu6 & Miniu6);
assign Ckniu6 = (Pgniu6 & Ajniu6);
assign Pgniu6 = (!Tiniu6);
assign Fhphu6 = (Ickiu6 ? vis_r2_o[28] : Gfniu6);
assign Ickiu6 = (~(Miniu6 & Jkniu6));
assign Miniu6 = (~(Ojniu6 | Qkniu6));
assign Ygphu6 = (Gumiu6 ? Gfniu6 : vis_r1_o[28]);
assign Gumiu6 = (Llniu6 & Igniu6);
assign Igniu6 = (Qkniu6 & Ajniu6);
assign Llniu6 = (~(Ojniu6 | Tiniu6));
assign Rgphu6 = (Numiu6 ? Gfniu6 : vis_r0_o[28]);
assign Numiu6 = (Slniu6 & Qkniu6);
assign Qkniu6 = (!Yhniu6);
assign Yhniu6 = (Zlniu6 | Gmniu6);
assign Zlniu6 = (~(HREADY & Nmniu6));
assign Slniu6 = (Wgniu6 & Jkniu6);
assign Jkniu6 = (~(Ajniu6 | Tiniu6));
assign Tiniu6 = (~(Umniu6 & Bnniu6));
assign Bnniu6 = (Inniu6 & Pnniu6);
assign Pnniu6 = (~(S8fpw6[10] & Wnniu6));
assign Inniu6 = (Doniu6 & Koniu6);
assign Koniu6 = (Roniu6 | Yoniu6);
assign Doniu6 = (Fpniu6 | Mpniu6);
assign Ajniu6 = (~(Tpniu6 & Aqniu6));
assign Aqniu6 = (Hqniu6 & Oqniu6);
assign Oqniu6 = (Vqniu6 | Mpniu6);
assign Hqniu6 = (~(S8fpw6[8] & Wnniu6));
assign Tpniu6 = (Crniu6 & Jrniu6);
assign Jrniu6 = (Qrniu6 | Yoniu6);
assign Wgniu6 = (!Ojniu6);
assign Ojniu6 = (~(Umniu6 & Xrniu6));
assign Xrniu6 = (Esniu6 & Lsniu6);
assign Lsniu6 = (Ssniu6 | Mpniu6);
assign Esniu6 = (Zsniu6 & Gtniu6);
assign Gtniu6 = (~(S8fpw6[11] & Wnniu6));
assign Zsniu6 = (Ntniu6 | Yoniu6);
assign Umniu6 = (Crniu6 & Utniu6);
assign Crniu6 = (Buniu6 & HREADY);
assign Buniu6 = (Nmniu6 & Iuniu6);
assign Nmniu6 = (~(Puniu6 & Wuniu6));
assign Wuniu6 = (Dvniu6 & Kvniu6);
assign Kvniu6 = (Rvniu6 & Yvniu6);
assign Yvniu6 = (~(Fwniu6 & Toaiu6));
assign Fwniu6 = (~(Knaiu6 | Cyfpw6[4]));
assign Rvniu6 = (Mwniu6 & Twniu6);
assign Dvniu6 = (Axniu6 & Hxniu6);
assign Hxniu6 = (~(Oxniu6 & Vxniu6));
assign Axniu6 = (Cyniu6 & Jyniu6);
assign Jyniu6 = (~(Qyniu6 & Xyniu6));
assign Xyniu6 = (~(Ezniu6 & Lzniu6));
assign Lzniu6 = (Szniu6 | Nlaiu6);
assign Cyniu6 = (~(Zzniu6 & Pugiu6));
assign Puniu6 = (G0oiu6 & N0oiu6);
assign N0oiu6 = (U0oiu6 & B1oiu6);
assign B1oiu6 = (~(Y0jiu6 & Wp0iu6));
assign U0oiu6 = (I1oiu6 & P1oiu6);
assign P1oiu6 = (~(W1oiu6 & Geaiu6));
assign W1oiu6 = (~(D2oiu6 & K2oiu6));
assign K2oiu6 = (~(R2oiu6 & Fd0iu6));
assign R2oiu6 = (~(Y2oiu6 | Knaiu6));
assign D2oiu6 = (F3oiu6 & M3oiu6);
assign M3oiu6 = (~(T3oiu6 & Md0iu6));
assign T3oiu6 = (~(A4oiu6 | Y7ghu6));
assign F3oiu6 = (~(H4oiu6 & O4oiu6));
assign I1oiu6 = (~(Imaiu6 & V4oiu6));
assign V4oiu6 = (~(C5oiu6 & J5oiu6));
assign J5oiu6 = (Q5oiu6 & X5oiu6);
assign Q5oiu6 = (~(E6oiu6 & Cyfpw6[4]));
assign C5oiu6 = (L6oiu6 & S6oiu6);
assign S6oiu6 = (~(Pthiu6 & Cyfpw6[7]));
assign L6oiu6 = (Tr0iu6 ? G7oiu6 : Z6oiu6);
assign G0oiu6 = (N7oiu6 & U7oiu6);
assign U7oiu6 = (Cyfpw6[6] ? I8oiu6 : B8oiu6);
assign I8oiu6 = (~(P8oiu6 & Zraiu6));
assign B8oiu6 = (W8oiu6 | D9oiu6);
assign N7oiu6 = (K9oiu6 & R9oiu6);
assign R9oiu6 = (~(Pthiu6 & Mfjiu6));
assign K9oiu6 = (H4ghu6 ? Faoiu6 : Y9oiu6);
assign Faoiu6 = (Maoiu6 & Taoiu6);
assign Taoiu6 = (~(Whfiu6 & Pthiu6));
assign Maoiu6 = (Aboiu6 & Hboiu6);
assign Hboiu6 = (~(Oboiu6 & Vboiu6));
assign Oboiu6 = (~(Ccoiu6 | Qxaiu6));
assign Aboiu6 = (~(Pugiu6 & Jcoiu6));
assign Jcoiu6 = (~(Qcoiu6 & Xcoiu6));
assign Xcoiu6 = (~(Edoiu6 & Ldoiu6));
assign Edoiu6 = (~(Jcaiu6 | Ii0iu6));
assign Y9oiu6 = (Sdoiu6 & Zdoiu6);
assign Zdoiu6 = (~(Geoiu6 & Neoiu6));
assign Sdoiu6 = (Ueoiu6 & Bfoiu6);
assign Bfoiu6 = (~(Ifoiu6 & Pfoiu6));
assign Ifoiu6 = (~(Wfoiu6 | Y7ghu6));
assign Ueoiu6 = (~(Dgoiu6 & Fd0iu6));
assign Dgoiu6 = (~(Ezniu6 | Cyfpw6[4]));
assign Gfniu6 = (~(Acniu6 & Kgoiu6));
assign Kgphu6 = (Y5liu6 ? Rgoiu6 : vis_apsr_o[3]);
assign Y5liu6 = (HREADY & Ygoiu6);
assign Ygoiu6 = (~(Fhoiu6 & Ug8iu6));
assign Rgoiu6 = (~(Mhoiu6 & Thoiu6));
assign Thoiu6 = (~(Ph8iu6 & Aioiu6));
assign Mhoiu6 = (Hioiu6 & Oioiu6);
assign Oioiu6 = (O7liu6 | Vioiu6);
assign O7liu6 = (!Ug8iu6);
assign Ug8iu6 = (~(Ph8iu6 | Yi8iu6));
assign Yi8iu6 = (!Cs8iu6);
assign Ph8iu6 = (!Hcniu6);
assign Hcniu6 = (Cjoiu6 & Vr8iu6);
assign Vr8iu6 = (~(Jjoiu6 & Wofiu6));
assign Cjoiu6 = (~(Jjoiu6 & Qjoiu6));
assign Hioiu6 = (Cs8iu6 | Ualiu6);
assign Cs8iu6 = (Mjfiu6 | Uzaiu6);
assign Uzaiu6 = (Xjoiu6 & Ekoiu6);
assign Ekoiu6 = (Lkoiu6 & Skoiu6);
assign Skoiu6 = (~(Zkoiu6 & Gloiu6));
assign Gloiu6 = (~(Nloiu6 | Xe8iu6));
assign Zkoiu6 = (~(G7oiu6 | Zraiu6));
assign Lkoiu6 = (Twniu6 & Uloiu6);
assign Xjoiu6 = (Bmoiu6 & Imoiu6);
assign Bmoiu6 = (~(L0niu6 & Tfjiu6));
assign Dgphu6 = (~(Pmoiu6 & Wmoiu6));
assign Wmoiu6 = (Dnoiu6 & Knoiu6);
assign Knoiu6 = (~(Ok8iu6 & vis_pc_o[30]));
assign Ok8iu6 = (Rnoiu6 & W8aiu6);
assign Rnoiu6 = (Ynoiu6 & Lm8iu6);
assign Ynoiu6 = (~(Fooiu6 & Lraiu6));
assign Fooiu6 = (Mooiu6 & Tr0iu6);
assign Mooiu6 = (Ttciu6 | D7fpw6[3]);
assign Dnoiu6 = (Tooiu6 & Apoiu6);
assign Apoiu6 = (~(Jl8iu6 & Ef1iu6));
assign Jl8iu6 = (Hpoiu6 & Lm8iu6);
assign Hpoiu6 = (~(Y7ghu6 & Opoiu6));
assign Opoiu6 = (Jojiu6 | Cyfpw6[1]);
assign Tooiu6 = (~(vis_apsr_o[3] & Ql8iu6));
assign Ql8iu6 = (Vpoiu6 & U19iu6);
assign U19iu6 = (Cqoiu6 & Jqoiu6);
assign Jqoiu6 = (~(Qqoiu6 & Xqoiu6));
assign Xqoiu6 = (~(V4aiu6 | R2aiu6));
assign Qqoiu6 = (~(Q5aiu6 | Prjiu6));
assign Cqoiu6 = (Eroiu6 & Lroiu6);
assign Eroiu6 = (~(Sroiu6 & Zroiu6));
assign Sroiu6 = (D7fpw6[8] & Nbkiu6);
assign Vpoiu6 = (Frliu6 & Lm8iu6);
assign Frliu6 = (~(Twniu6 & Gsoiu6));
assign Gsoiu6 = (~(Nsoiu6 & Usoiu6));
assign Usoiu6 = (Btoiu6 & D7fpw6[3]);
assign Nsoiu6 = (~(Q5aiu6 | Ttciu6));
assign Pmoiu6 = (Itoiu6 & Ptoiu6);
assign Ptoiu6 = (Lm8iu6 | Wtoiu6);
assign Lm8iu6 = (!W29iu6);
assign W29iu6 = (Duoiu6 & Hx9iu6);
assign Duoiu6 = (~(HREADY & Kuoiu6));
assign Kuoiu6 = (~(Ruoiu6 & Yuoiu6));
assign Yuoiu6 = (Fvoiu6 & Mvoiu6);
assign Mvoiu6 = (Tvoiu6 & Awoiu6);
assign Awoiu6 = (~(Hwoiu6 & Ia8iu6));
assign Hwoiu6 = (Vviiu6 & D7fpw6[12]);
assign Tvoiu6 = (~(Y0jiu6 & Owoiu6));
assign Fvoiu6 = (Vwoiu6 & Cxoiu6);
assign Cxoiu6 = (Jxoiu6 | Qxoiu6);
assign Vwoiu6 = (~(Xxoiu6 & Zraiu6));
assign Xxoiu6 = (~(Eyoiu6 & Lyoiu6));
assign Lyoiu6 = (Syoiu6 & Td0iu6);
assign Syoiu6 = (~(Zyoiu6 & Gzoiu6));
assign Gzoiu6 = (~(Lraiu6 | Nzoiu6));
assign Zyoiu6 = (Wliiu6 & Dmiiu6);
assign Eyoiu6 = (Uzoiu6 & B0piu6);
assign B0piu6 = (~(I0piu6 & P0piu6));
assign I0piu6 = (W0piu6 & D7fpw6[13]);
assign Uzoiu6 = (~(Vxniu6 & D1piu6));
assign Ruoiu6 = (K1piu6 & R1piu6);
assign R1piu6 = (Y1piu6 & F2piu6);
assign F2piu6 = (~(L0niu6 & M2piu6));
assign L0niu6 = (T2piu6 & Md0iu6);
assign T2piu6 = (~(A4oiu6 | Mr0iu6));
assign Y1piu6 = (~(Geoiu6 & Qe8iu6));
assign K1piu6 = (A3piu6 & F85iu6);
assign A3piu6 = (Cyfpw6[3] ? O3piu6 : H3piu6);
assign O3piu6 = (~(V3piu6 & W8aiu6));
assign V3piu6 = (C4piu6 & Nlaiu6);
assign C4piu6 = (~(Lraiu6 & J4piu6));
assign J4piu6 = (~(Q4piu6 & T0hhu6));
assign Q4piu6 = (X4piu6 & Ftjiu6);
assign X4piu6 = (V4aiu6 | R9aiu6);
assign Itoiu6 = (~(Zm8iu6 & Lm1iu6));
assign Zm8iu6 = (!Hx9iu6);
assign Hx9iu6 = (~(E5piu6 & HALTED));
assign E5piu6 = (Ar1iu6 & Npdhu6);
assign Wfphu6 = (L5piu6 | Ln7iu6);
assign L5piu6 = (Zn7iu6 ? T15iu6 : Ppfpw6[16]);
assign Zn7iu6 = (~(A2ciu6 & S5piu6));
assign S5piu6 = (~(Z5piu6 & G6piu6));
assign G6piu6 = (~(N6piu6 | C0ehu6));
assign Z5piu6 = (~(Qqhiu6 | Juzhu6));
assign A2ciu6 = (!Ln7iu6);
assign Ln7iu6 = (H2ciu6 | Ivfhu6);
assign H2ciu6 = (!Jm7iu6);
assign Jm7iu6 = (Wofiu6 | U6piu6);
assign T15iu6 = (~(Svdpw6 & Vobiu6));
assign Pfphu6 = (Ex4iu6 | B7piu6);
assign B7piu6 = (Dhgpw6[0] & I7piu6);
assign I7piu6 = (~(Scbiu6 & T24iu6));
assign Ex4iu6 = (~(P7piu6 & W7piu6));
assign W7piu6 = (~(D8piu6 & Tu4iu6));
assign Tu4iu6 = (K8piu6 & R8piu6);
assign R8piu6 = (Y8piu6 & F9piu6);
assign F9piu6 = (M9piu6 & T9piu6);
assign T9piu6 = (Aapiu6 & Asliu6);
assign Aapiu6 = (~(W74iu6 | I74iu6));
assign M9piu6 = (~(Y84iu6 | R84iu6));
assign Y8piu6 = (Hapiu6 & Oapiu6);
assign Oapiu6 = (~(T94iu6 | F94iu6));
assign Hapiu6 = (Lm1iu6 & Rykiu6);
assign K8piu6 = (Vapiu6 & Cbpiu6);
assign Cbpiu6 = (Jbpiu6 & Qbpiu6);
assign Qbpiu6 = (Xbpiu6 & P74iu6);
assign Xbpiu6 = (M94iu6 & Z54iu6);
assign Jbpiu6 = (U64iu6 & B74iu6);
assign Vapiu6 = (Ecpiu6 & Lcpiu6);
assign Lcpiu6 = (G64iu6 & N64iu6);
assign Ecpiu6 = (~(Duhiu6 | Ps4iu6));
assign D8piu6 = (T24iu6 & O34iu6);
assign P7piu6 = (~(Scpiu6 & Zcpiu6));
assign Zcpiu6 = (Gdpiu6 & Jehhu6);
assign Gdpiu6 = (Ndpiu6 & Udpiu6);
assign Ndpiu6 = (~(Bepiu6 & Zrhiu6));
assign Zrhiu6 = (~(LOCKUP | C0ehu6));
assign Bepiu6 = (Uc5iu6 & Sb5iu6);
assign Uc5iu6 = (~(Iepiu6 & K2aiu6));
assign Scpiu6 = (Hbhhu6 & HREADY);
assign Ifphu6 = (~(Pepiu6 & Wepiu6));
assign Wepiu6 = (~(Dfpiu6 & Lx4iu6));
assign Lx4iu6 = (Kfpiu6 | Rfpiu6);
assign Dfpiu6 = (~(Eh6iu6 & Yfpiu6));
assign Pepiu6 = (~(Dhgpw6[2] & Yfpiu6));
assign Yfpiu6 = (~(Scbiu6 & Ud4iu6));
assign Scbiu6 = (Fgpiu6 & A2nhu6);
assign Bfphu6 = (~(Mgpiu6 & Tgpiu6));
assign Tgpiu6 = (~(Rfpiu6 & Ahpiu6));
assign Ahpiu6 = (~(Eh6iu6 & Hhpiu6));
assign Rfpiu6 = (Ohpiu6 & Yuhhu6);
assign Ohpiu6 = (~(E81iu6 | Vhpiu6));
assign Vhpiu6 = (Cipiu6 & Jipiu6);
assign Jipiu6 = (~(Qipiu6 & Xipiu6));
assign Qipiu6 = (Ejpiu6 ? Lwgpw6[0] : Lwgpw6[1]);
assign Cipiu6 = (Ljpiu6 | Ty0iu6);
assign Ty0iu6 = (Lwgpw6[0] | Lwgpw6[1]);
assign E81iu6 = (~(Sjpiu6 & Lwgpw6[2]));
assign Mgpiu6 = (~(Hwmhu6 & Hhpiu6));
assign Hhpiu6 = (~(Ws4iu6 & Ps4iu6));
assign Uephu6 = (~(Zjpiu6 & Gkpiu6));
assign Gkpiu6 = (~(Kfpiu6 & Nkpiu6));
assign Nkpiu6 = (~(Eh6iu6 & Ukpiu6));
assign Kfpiu6 = (Blpiu6 & Mekhu6);
assign Blpiu6 = (~(Yx0iu6 | Ilpiu6));
assign Ilpiu6 = (Plpiu6 & Wlpiu6);
assign Wlpiu6 = (~(Dmpiu6 & Xipiu6));
assign Xipiu6 = (Kmpiu6 & Rmpiu6);
assign Rmpiu6 = (Z18iu6 | Ympiu6);
assign Kmpiu6 = (~(HMASTER | L18iu6));
assign Dmpiu6 = (Fnpiu6 ? R2hpw6[1] : R2hpw6[0]);
assign Plpiu6 = (Ljpiu6 | Nv0iu6);
assign Nv0iu6 = (R2hpw6[0] | R2hpw6[1]);
assign Ljpiu6 = (~(Mnpiu6 & Sufpw6[1]));
assign Mnpiu6 = (Sufpw6[0] & K9aiu6);
assign Yx0iu6 = (~(Sjpiu6 & R2hpw6[2]));
assign Sjpiu6 = (E5hhu6 & Jehhu6);
assign Zjpiu6 = (~(Vxmhu6 & Ukpiu6));
assign Ukpiu6 = (~(Eg7iu6 & Ps4iu6));
assign Ps4iu6 = (!A2nhu6);
assign Nephu6 = (~(Tnpiu6 & Aopiu6));
assign Aopiu6 = (Hopiu6 & Oopiu6);
assign Oopiu6 = (~(Tnhpw6[1] & Bo1iu6));
assign Hopiu6 = (Vopiu6 & Po1iu6);
assign Vopiu6 = (~(Wo1iu6 & Cppiu6));
assign Cppiu6 = (~(Jppiu6 & Qppiu6));
assign Qppiu6 = (Xppiu6 & Eqpiu6);
assign Eqpiu6 = (Lqpiu6 & Sqpiu6);
assign Sqpiu6 = (Zqpiu6 & Grpiu6);
assign Grpiu6 = (~(R2hpw6[1] & Eg7iu6));
assign Zqpiu6 = (~(Dhgpw6[1] & Fgpiu6));
assign Lqpiu6 = (Nrpiu6 & Urpiu6);
assign Urpiu6 = (~(G4hpw6[1] & Sg7iu6));
assign Nrpiu6 = (~(Aygpw6[1] & Jf7iu6));
assign Xppiu6 = (Bspiu6 & Ispiu6);
assign Ispiu6 = (~(Ar1iu6 & Fkfpw6[1]));
assign Bspiu6 = (Pspiu6 & Wspiu6);
assign Wspiu6 = (Duhiu6 | Udpiu6);
assign Pspiu6 = (~(Lwgpw6[1] & Ws4iu6));
assign Jppiu6 = (Dtpiu6 & Ktpiu6);
assign Ktpiu6 = (Rtpiu6 & Ytpiu6);
assign Ytpiu6 = (Fupiu6 & Mupiu6);
assign Mupiu6 = (~(HRDATA[1] & St1iu6));
assign Fupiu6 = (~(Zt1iu6 & Pzgpw6[1]));
assign Rtpiu6 = (Tupiu6 & Avpiu6);
assign Avpiu6 = (~(Kw1iu6 & V5hpw6[1]));
assign Tupiu6 = (~(Iv1iu6 & vis_pc_o[0]));
assign Dtpiu6 = (Hvpiu6 & Ovpiu6);
assign Hvpiu6 = (Vvpiu6 & Yw1iu6);
assign Tnpiu6 = (Cwpiu6 & Jwpiu6);
assign Jwpiu6 = (~(Qwpiu6 & Aphpw6[2]));
assign Cwpiu6 = (~(Uthpw6[1] & Sf1iu6));
assign Gephu6 = (~(Xwpiu6 & Expiu6));
assign Expiu6 = (~(Uthpw6[2] & Sf1iu6));
assign Xwpiu6 = (Lxpiu6 & Sxpiu6);
assign Sxpiu6 = (~(Wo1iu6 & Zxpiu6));
assign Zxpiu6 = (~(Gypiu6 & Nypiu6));
assign Nypiu6 = (Uypiu6 & Bzpiu6);
assign Bzpiu6 = (Izpiu6 & Pzpiu6);
assign Pzpiu6 = (Wzpiu6 & D0qiu6);
assign D0qiu6 = (~(K0qiu6 & Hbhhu6));
assign K0qiu6 = (~(Duhiu6 | Zwciu6));
assign Izpiu6 = (R0qiu6 & Y0qiu6);
assign Y0qiu6 = (~(Eg7iu6 & R2hpw6[2]));
assign R0qiu6 = (F1qiu6 & M1qiu6);
assign M1qiu6 = (~(T1qiu6 & A2qiu6));
assign T1qiu6 = (X8hpw6[5] ? O2qiu6 : H2qiu6);
assign O2qiu6 = (V2qiu6 | C3qiu6);
assign V2qiu6 = (Dr6iu6 & Vm6iu6);
assign H2qiu6 = (~(J3qiu6 | Dr6iu6));
assign F1qiu6 = (~(Q3qiu6 & Fl6iu6));
assign Uypiu6 = (X3qiu6 & E4qiu6);
assign E4qiu6 = (L4qiu6 & S4qiu6);
assign S4qiu6 = (~(Aygpw6[2] & Jf7iu6));
assign L4qiu6 = (Z4qiu6 & G5qiu6);
assign G5qiu6 = (~(Dhgpw6[2] & Fgpiu6));
assign Z4qiu6 = (~(G4hpw6[2] & Sg7iu6));
assign X3qiu6 = (N5qiu6 & U5qiu6);
assign U5qiu6 = (~(Togpw6[2] & Vr1iu6));
assign N5qiu6 = (~(Ws4iu6 & Lwgpw6[2]));
assign Gypiu6 = (B6qiu6 & I6qiu6);
assign I6qiu6 = (P6qiu6 & W6qiu6);
assign W6qiu6 = (D7qiu6 & K7qiu6);
assign K7qiu6 = (~(HRDATA[2] & St1iu6));
assign D7qiu6 = (R7qiu6 & Y7qiu6);
assign Y7qiu6 = (~(Gtgpw6[2] & Cs1iu6));
assign R7qiu6 = (~(Ar1iu6 & Fkfpw6[2]));
assign P6qiu6 = (F8qiu6 & M8qiu6);
assign M8qiu6 = (~(E1hpw6[2] & Zt1iu6));
assign F8qiu6 = (~(Gqgpw6[2] & Xs1iu6));
assign B6qiu6 = (T8qiu6 & A9qiu6);
assign A9qiu6 = (H9qiu6 & O9qiu6);
assign O9qiu6 = (~(Iv1iu6 & vis_pc_o[1]));
assign H9qiu6 = (V9qiu6 & Caqiu6);
assign Caqiu6 = (~(Trgpw6[2] & Dw1iu6));
assign V9qiu6 = (~(K7hpw6[2] & Kw1iu6));
assign T8qiu6 = (Jaqiu6 & Qaqiu6);
assign Lxpiu6 = (~(Tnhpw6[2] & Bo1iu6));
assign Zdphu6 = (~(Xaqiu6 & Ebqiu6));
assign Ebqiu6 = (~(Uthpw6[3] & Sf1iu6));
assign Xaqiu6 = (Lbqiu6 & Sbqiu6);
assign Sbqiu6 = (~(Wo1iu6 & Zbqiu6));
assign Zbqiu6 = (~(Gcqiu6 & Ncqiu6));
assign Ncqiu6 = (Ucqiu6 & Bdqiu6);
assign Bdqiu6 = (Idqiu6 & Pdqiu6);
assign Pdqiu6 = (Wdqiu6 & Deqiu6);
assign Deqiu6 = (~(Dhgpw6[3] & Fgpiu6));
assign Wdqiu6 = (Keqiu6 & Reqiu6);
assign Keqiu6 = (~(Yeqiu6 & Ffqiu6));
assign Yeqiu6 = (~(Mfqiu6 | X8hpw6[0]));
assign Idqiu6 = (Tfqiu6 & Agqiu6);
assign Agqiu6 = (~(G4hpw6[3] & Sg7iu6));
assign Tfqiu6 = (~(Aygpw6[3] & Jf7iu6));
assign Ucqiu6 = (Hgqiu6 & Ogqiu6);
assign Ogqiu6 = (Vgqiu6 & Chqiu6);
assign Chqiu6 = (~(Togpw6[3] & Vr1iu6));
assign Vgqiu6 = (Jhqiu6 | Duhiu6);
assign Hgqiu6 = (Qhqiu6 & Xhqiu6);
assign Xhqiu6 = (~(Gtgpw6[3] & Cs1iu6));
assign Qhqiu6 = (~(Ar1iu6 & Fkfpw6[3]));
assign Gcqiu6 = (Eiqiu6 & Liqiu6);
assign Liqiu6 = (Siqiu6 & Ziqiu6);
assign Ziqiu6 = (Gjqiu6 & Njqiu6);
assign Njqiu6 = (~(Gqgpw6[3] & Xs1iu6));
assign Gjqiu6 = (Ujqiu6 & Bkqiu6);
assign Bkqiu6 = (~(HRDATA[3] & St1iu6));
assign Ujqiu6 = (~(E1hpw6[3] & Zt1iu6));
assign Siqiu6 = (Ikqiu6 & Pkqiu6);
assign Pkqiu6 = (~(Trgpw6[3] & Dw1iu6));
assign Ikqiu6 = (~(K7hpw6[3] & Kw1iu6));
assign Eiqiu6 = (Wkqiu6 & Dlqiu6);
assign Dlqiu6 = (Vvpiu6 & Klqiu6);
assign Klqiu6 = (~(Iv1iu6 & vis_pc_o[2]));
assign Vvpiu6 = (~(Rlqiu6 | Ylqiu6));
assign Rlqiu6 = (X8hpw6[4] ? Q3qiu6 : Fmqiu6);
assign Fmqiu6 = (Mmqiu6 & X8hpw6[1]);
assign Wkqiu6 = (Tmqiu6 & Anqiu6);
assign Lbqiu6 = (~(Tnhpw6[3] & Bo1iu6));
assign Sdphu6 = (~(Hnqiu6 & Onqiu6));
assign Onqiu6 = (Vnqiu6 & Coqiu6);
assign Coqiu6 = (~(Wo1iu6 & Joqiu6));
assign Joqiu6 = (~(Qoqiu6 & Xoqiu6));
assign Xoqiu6 = (Epqiu6 & Lpqiu6);
assign Lpqiu6 = (Spqiu6 & Zpqiu6);
assign Zpqiu6 = (Gqqiu6 & Nqqiu6);
assign Nqqiu6 = (~(ECOREVNUM[16] & Uqqiu6));
assign Gqqiu6 = (Brqiu6 & Irqiu6);
assign Brqiu6 = (~(ECOREVNUM[12] & Prqiu6));
assign Spqiu6 = (Wrqiu6 & Dsqiu6);
assign Dsqiu6 = (~(ECOREVNUM[4] & Ksqiu6));
assign Wrqiu6 = (~(ECOREVNUM[8] & Rsqiu6));
assign Epqiu6 = (Ysqiu6 & Ftqiu6);
assign Ftqiu6 = (Mtqiu6 & Ttqiu6);
assign Ttqiu6 = (~(Aygpw6[4] & Jf7iu6));
assign Mtqiu6 = (Auqiu6 & Huqiu6);
assign Huqiu6 = (~(Dhgpw6[4] & Fgpiu6));
assign Auqiu6 = (~(G4hpw6[4] & Sg7iu6));
assign Ysqiu6 = (Ouqiu6 & Vuqiu6);
assign Vuqiu6 = (~(Togpw6[4] & Vr1iu6));
assign Ouqiu6 = (~(Gtgpw6[4] & Cs1iu6));
assign Qoqiu6 = (Cvqiu6 & Jvqiu6);
assign Jvqiu6 = (Qvqiu6 & Xvqiu6);
assign Xvqiu6 = (Ewqiu6 & Lwqiu6);
assign Lwqiu6 = (~(E1hpw6[4] & Zt1iu6));
assign Ewqiu6 = (Swqiu6 & Zwqiu6);
assign Zwqiu6 = (~(Ar1iu6 & Fkfpw6[4]));
assign Swqiu6 = (~(HRDATA[4] & St1iu6));
assign Qvqiu6 = (Gxqiu6 & Nxqiu6);
assign Nxqiu6 = (~(Gqgpw6[4] & Xs1iu6));
assign Gxqiu6 = (~(Trgpw6[4] & Dw1iu6));
assign Cvqiu6 = (Uxqiu6 & Byqiu6);
assign Byqiu6 = (Iyqiu6 & Pyqiu6);
assign Pyqiu6 = (~(Wyqiu6 & Dzqiu6));
assign Iyqiu6 = (Kzqiu6 & Rzqiu6);
assign Rzqiu6 = (~(K7hpw6[4] & Kw1iu6));
assign Kzqiu6 = (~(vis_pc_o[3] & Iv1iu6));
assign Uxqiu6 = (Yzqiu6 & F0riu6);
assign Vnqiu6 = (~(Jshpw6[4] & Bo1iu6));
assign Hnqiu6 = (M0riu6 & T0riu6);
assign T0riu6 = (~(Qwpiu6 & Cynhu6));
assign M0riu6 = (~(Uthpw6[4] & Sf1iu6));
assign Ldphu6 = (~(A1riu6 & H1riu6));
assign H1riu6 = (O1riu6 & V1riu6);
assign O1riu6 = (~(Wo1iu6 & C2riu6));
assign C2riu6 = (~(J2riu6 & Q2riu6));
assign Q2riu6 = (X2riu6 & E3riu6);
assign E3riu6 = (L3riu6 & S3riu6);
assign S3riu6 = (Z3riu6 & G4riu6);
assign G4riu6 = (~(ECOREVNUM[17] & Uqqiu6));
assign Z3riu6 = (N4riu6 & Irqiu6);
assign Irqiu6 = (!U4riu6);
assign N4riu6 = (~(ECOREVNUM[13] & Prqiu6));
assign L3riu6 = (B5riu6 & I5riu6);
assign I5riu6 = (~(ECOREVNUM[5] & Ksqiu6));
assign B5riu6 = (~(ECOREVNUM[9] & Rsqiu6));
assign X2riu6 = (P5riu6 & W5riu6);
assign W5riu6 = (D6riu6 & K6riu6);
assign K6riu6 = (~(Togpw6[5] & Vr1iu6));
assign D6riu6 = (~(Gtgpw6[5] & Cs1iu6));
assign P5riu6 = (R6riu6 & Y6riu6);
assign Y6riu6 = (~(Ar1iu6 & Fkfpw6[5]));
assign R6riu6 = (~(HRDATA[5] & St1iu6));
assign J2riu6 = (F7riu6 & M7riu6);
assign M7riu6 = (T7riu6 & A8riu6);
assign A8riu6 = (H8riu6 & O8riu6);
assign O8riu6 = (~(E1hpw6[5] & Zt1iu6));
assign H8riu6 = (~(Gqgpw6[5] & Xs1iu6));
assign T7riu6 = (V8riu6 & C9riu6);
assign C9riu6 = (~(Trgpw6[5] & Dw1iu6));
assign V8riu6 = (~(K7hpw6[5] & Kw1iu6));
assign F7riu6 = (J9riu6 & Q9riu6);
assign Q9riu6 = (F0riu6 & X9riu6);
assign X9riu6 = (~(vis_pc_o[4] & Iv1iu6));
assign J9riu6 = (Eariu6 & Lariu6);
assign A1riu6 = (Sariu6 & Zariu6);
assign Zariu6 = (~(Jshpw6[5] & Bo1iu6));
assign Sariu6 = (~(Uthpw6[5] & Sf1iu6));
assign Edphu6 = (~(Gbriu6 & Nbriu6));
assign Nbriu6 = (Ubriu6 & Bcriu6);
assign Ubriu6 = (~(Wo1iu6 & Icriu6));
assign Icriu6 = (~(Pcriu6 & Wcriu6));
assign Wcriu6 = (Ddriu6 & Kdriu6);
assign Kdriu6 = (Rdriu6 & Ydriu6);
assign Ydriu6 = (Feriu6 & Reqiu6);
assign Feriu6 = (~(U4riu6 | Ve7iu6));
assign Rdriu6 = (Meriu6 & Teriu6);
assign Teriu6 = (~(ECOREVNUM[14] & Prqiu6));
assign Meriu6 = (~(ECOREVNUM[18] & Uqqiu6));
assign Ddriu6 = (Afriu6 & Hfriu6);
assign Hfriu6 = (Ofriu6 & Vfriu6);
assign Vfriu6 = (~(ECOREVNUM[6] & Ksqiu6));
assign Ofriu6 = (~(ECOREVNUM[10] & Rsqiu6));
assign Afriu6 = (Cgriu6 & Jgriu6);
assign Jgriu6 = (~(Togpw6[6] & Vr1iu6));
assign Cgriu6 = (~(Gtgpw6[6] & Cs1iu6));
assign Pcriu6 = (Qgriu6 & Xgriu6);
assign Xgriu6 = (Ehriu6 & Lhriu6);
assign Lhriu6 = (Shriu6 & Zhriu6);
assign Zhriu6 = (~(E1hpw6[6] & Zt1iu6));
assign Shriu6 = (Giriu6 & Niriu6);
assign Niriu6 = (~(Ar1iu6 & Fkfpw6[6]));
assign Giriu6 = (~(HRDATA[6] & St1iu6));
assign Ehriu6 = (Uiriu6 & Bjriu6);
assign Bjriu6 = (~(Gqgpw6[6] & Xs1iu6));
assign Uiriu6 = (~(Trgpw6[6] & Dw1iu6));
assign Qgriu6 = (Ijriu6 & Pjriu6);
assign Pjriu6 = (Wjriu6 & Dkriu6);
assign Dkriu6 = (~(K7hpw6[6] & Kw1iu6));
assign Wjriu6 = (~(vis_pc_o[5] & Iv1iu6));
assign Ijriu6 = (Kkriu6 & Lariu6);
assign Gbriu6 = (Rkriu6 & Ykriu6);
assign Ykriu6 = (~(Jshpw6[6] & Bo1iu6));
assign Rkriu6 = (~(Uthpw6[6] & Sf1iu6));
assign Xcphu6 = (~(Flriu6 & Mlriu6));
assign Mlriu6 = (~(Uthpw6[7] & Sf1iu6));
assign Flriu6 = (Tlriu6 & Amriu6);
assign Amriu6 = (~(Wo1iu6 & Hmriu6));
assign Hmriu6 = (~(Omriu6 & Vmriu6));
assign Vmriu6 = (Cnriu6 & Jnriu6);
assign Jnriu6 = (Qnriu6 & Xnriu6);
assign Xnriu6 = (Eoriu6 & Loriu6);
assign Loriu6 = (~(ECOREVNUM[15] & Prqiu6));
assign Prqiu6 = (Soriu6 & A2qiu6);
assign Soriu6 = (Dzqiu6 & Cvciu6);
assign Eoriu6 = (~(ECOREVNUM[19] & Uqqiu6));
assign Uqqiu6 = (Zoriu6 & Wyqiu6);
assign Zoriu6 = (~(Fl6iu6 | Mfqiu6));
assign Qnriu6 = (Gpriu6 & Npriu6);
assign Npriu6 = (~(ECOREVNUM[7] & Ksqiu6));
assign Ksqiu6 = (Upriu6 & A2qiu6);
assign Upriu6 = (Bqriu6 & Cvciu6);
assign Gpriu6 = (~(ECOREVNUM[11] & Rsqiu6));
assign Rsqiu6 = (Iqriu6 & X8hpw6[4]);
assign Cnriu6 = (Pqriu6 & Wqriu6);
assign Wqriu6 = (Drriu6 & Krriu6);
assign Krriu6 = (~(Togpw6[7] & Vr1iu6));
assign Drriu6 = (~(Gtgpw6[7] & Cs1iu6));
assign Pqriu6 = (Rrriu6 & Yrriu6);
assign Yrriu6 = (~(Ar1iu6 & Fkfpw6[7]));
assign Rrriu6 = (~(HRDATA[7] & St1iu6));
assign Omriu6 = (Fsriu6 & Msriu6);
assign Msriu6 = (Tsriu6 & Atriu6);
assign Atriu6 = (Htriu6 & Otriu6);
assign Otriu6 = (~(E1hpw6[7] & Zt1iu6));
assign Htriu6 = (~(Gqgpw6[7] & Xs1iu6));
assign Tsriu6 = (Vtriu6 & Curiu6);
assign Curiu6 = (~(Trgpw6[7] & Dw1iu6));
assign Vtriu6 = (~(K7hpw6[7] & Kw1iu6));
assign Fsriu6 = (Juriu6 & Quriu6);
assign Quriu6 = (F0riu6 & Xuriu6);
assign Xuriu6 = (~(vis_pc_o[6] & Iv1iu6));
assign F0riu6 = (Evriu6 & Lvriu6);
assign Lvriu6 = (Wzpiu6 & Svriu6);
assign Wzpiu6 = (Zvriu6 & Reqiu6);
assign Zvriu6 = (~(Gwriu6 & Wyqiu6));
assign Gwriu6 = (~(Nwriu6 | X8hpw6[4]));
assign Evriu6 = (Uwriu6 & Bxriu6);
assign Bxriu6 = (~(Ixriu6 & Fl6iu6));
assign Juriu6 = (Pxriu6 & Lariu6);
assign Lariu6 = (Wxriu6 & Dyriu6);
assign Dyriu6 = (~(Kyriu6 & Ixriu6));
assign Kyriu6 = (~(Fl6iu6 | Vm6iu6));
assign Wxriu6 = (~(Ryriu6 & Cvciu6));
assign Tlriu6 = (~(Jshpw6[7] & Bo1iu6));
assign Qcphu6 = (~(Yyriu6 & Fzriu6));
assign Fzriu6 = (~(Uthpw6[8] & Sf1iu6));
assign Yyriu6 = (Mzriu6 & Tzriu6);
assign Tzriu6 = (~(Wo1iu6 & A0siu6));
assign A0siu6 = (~(H0siu6 & O0siu6));
assign O0siu6 = (V0siu6 & C1siu6);
assign C1siu6 = (J1siu6 & Q1siu6);
assign Q1siu6 = (~(Gtgpw6[8] & Cs1iu6));
assign J1siu6 = (X1siu6 & Reqiu6);
assign X1siu6 = (~(Togpw6[8] & Vr1iu6));
assign V0siu6 = (E2siu6 & L2siu6);
assign L2siu6 = (~(E1hpw6[8] & Zt1iu6));
assign E2siu6 = (S2siu6 & Z2siu6);
assign Z2siu6 = (~(Ar1iu6 & Fkfpw6[8]));
assign S2siu6 = (~(HRDATA[8] & St1iu6));
assign H0siu6 = (G3siu6 & N3siu6);
assign N3siu6 = (U3siu6 & B4siu6);
assign B4siu6 = (~(K7hpw6[8] & Kw1iu6));
assign U3siu6 = (I4siu6 & P4siu6);
assign P4siu6 = (~(Gqgpw6[8] & Xs1iu6));
assign I4siu6 = (~(Trgpw6[8] & Dw1iu6));
assign G3siu6 = (W4siu6 & D5siu6);
assign D5siu6 = (~(vis_pc_o[7] & Iv1iu6));
assign Mzriu6 = (~(Jshpw6[8] & Bo1iu6));
assign Jcphu6 = (~(K5siu6 & R5siu6));
assign R5siu6 = (~(Uthpw6[9] & Sf1iu6));
assign K5siu6 = (Y5siu6 & F6siu6);
assign F6siu6 = (~(Wo1iu6 & M6siu6));
assign M6siu6 = (~(T6siu6 & A7siu6));
assign A7siu6 = (H7siu6 & O7siu6);
assign O7siu6 = (V7siu6 & C8siu6);
assign C8siu6 = (~(Gtgpw6[9] & Cs1iu6));
assign V7siu6 = (J8siu6 & Reqiu6);
assign J8siu6 = (~(Togpw6[9] & Vr1iu6));
assign H7siu6 = (Q8siu6 & X8siu6);
assign X8siu6 = (~(E1hpw6[9] & Zt1iu6));
assign Q8siu6 = (E9siu6 & L9siu6);
assign L9siu6 = (~(Ar1iu6 & Fkfpw6[9]));
assign E9siu6 = (~(HRDATA[9] & St1iu6));
assign T6siu6 = (S9siu6 & Z9siu6);
assign Z9siu6 = (Gasiu6 & Nasiu6);
assign Nasiu6 = (~(K7hpw6[9] & Kw1iu6));
assign Gasiu6 = (Uasiu6 & Bbsiu6);
assign Bbsiu6 = (~(Gqgpw6[9] & Xs1iu6));
assign Uasiu6 = (~(Trgpw6[9] & Dw1iu6));
assign S9siu6 = (Ibsiu6 & Pbsiu6);
assign Pbsiu6 = (~(vis_pc_o[8] & Iv1iu6));
assign Y5siu6 = (~(Jshpw6[9] & Bo1iu6));
assign Ccphu6 = (~(Wbsiu6 & Dcsiu6));
assign Dcsiu6 = (~(Uthpw6[10] & Sf1iu6));
assign Wbsiu6 = (Kcsiu6 & Rcsiu6);
assign Rcsiu6 = (~(Wo1iu6 & Ycsiu6));
assign Ycsiu6 = (~(Fdsiu6 & Mdsiu6));
assign Mdsiu6 = (Tdsiu6 & Aesiu6);
assign Aesiu6 = (Hesiu6 & Oesiu6);
assign Oesiu6 = (~(Togpw6[10] & Vr1iu6));
assign Hesiu6 = (Vesiu6 & Reqiu6);
assign Vesiu6 = (~(Yc7iu6 & S3hhu6));
assign Tdsiu6 = (Cfsiu6 & Jfsiu6);
assign Jfsiu6 = (~(HRDATA[10] & St1iu6));
assign Cfsiu6 = (Qfsiu6 & Xfsiu6);
assign Xfsiu6 = (~(Gtgpw6[10] & Cs1iu6));
assign Qfsiu6 = (~(Ar1iu6 & Fkfpw6[10]));
assign Fdsiu6 = (Egsiu6 & Lgsiu6);
assign Lgsiu6 = (Sgsiu6 & Zgsiu6);
assign Zgsiu6 = (~(Trgpw6[10] & Dw1iu6));
assign Sgsiu6 = (Ghsiu6 & Nhsiu6);
assign Nhsiu6 = (~(E1hpw6[10] & Zt1iu6));
assign Ghsiu6 = (~(Gqgpw6[10] & Xs1iu6));
assign Egsiu6 = (Uhsiu6 & Bisiu6);
assign Uhsiu6 = (Iisiu6 & Pisiu6);
assign Pisiu6 = (~(K7hpw6[10] & Kw1iu6));
assign Iisiu6 = (~(vis_pc_o[9] & Iv1iu6));
assign Kcsiu6 = (~(Jshpw6[10] & Bo1iu6));
assign Vbphu6 = (~(Wisiu6 & Djsiu6));
assign Djsiu6 = (~(Uthpw6[11] & Sf1iu6));
assign Wisiu6 = (Kjsiu6 & Rjsiu6);
assign Rjsiu6 = (~(Wo1iu6 & Yjsiu6));
assign Yjsiu6 = (~(Fksiu6 & Mksiu6));
assign Mksiu6 = (Tksiu6 & Alsiu6);
assign Alsiu6 = (Hlsiu6 & Olsiu6);
assign Olsiu6 = (~(Gtgpw6[11] & Cs1iu6));
assign Hlsiu6 = (Vlsiu6 & Reqiu6);
assign Vlsiu6 = (~(Togpw6[11] & Vr1iu6));
assign Tksiu6 = (Cmsiu6 & Jmsiu6);
assign Jmsiu6 = (~(E1hpw6[11] & Zt1iu6));
assign Cmsiu6 = (Qmsiu6 & Xmsiu6);
assign Xmsiu6 = (~(Ar1iu6 & Fkfpw6[11]));
assign Qmsiu6 = (~(HRDATA[11] & St1iu6));
assign Fksiu6 = (Ensiu6 & Lnsiu6);
assign Lnsiu6 = (Snsiu6 & Znsiu6);
assign Znsiu6 = (~(K7hpw6[11] & Kw1iu6));
assign Snsiu6 = (Gosiu6 & Nosiu6);
assign Nosiu6 = (~(Gqgpw6[11] & Xs1iu6));
assign Gosiu6 = (~(Trgpw6[11] & Dw1iu6));
assign Ensiu6 = (Uosiu6 & Bpsiu6);
assign Bpsiu6 = (~(vis_pc_o[10] & Iv1iu6));
assign Kjsiu6 = (~(Jshpw6[11] & Bo1iu6));
assign Obphu6 = (~(Ipsiu6 & Ppsiu6));
assign Ppsiu6 = (Wpsiu6 & Po1iu6);
assign Wpsiu6 = (~(Wo1iu6 & Dqsiu6));
assign Dqsiu6 = (~(Kqsiu6 & Rqsiu6));
assign Rqsiu6 = (Yqsiu6 & Frsiu6);
assign Frsiu6 = (Mrsiu6 & Trsiu6);
assign Trsiu6 = (~(Gtgpw6[12] & Cs1iu6));
assign Mrsiu6 = (Assiu6 & Hssiu6);
assign Assiu6 = (~(Togpw6[12] & Vr1iu6));
assign Yqsiu6 = (Ossiu6 & Vssiu6);
assign Vssiu6 = (~(E1hpw6[12] & Zt1iu6));
assign Ossiu6 = (Ctsiu6 & Jtsiu6);
assign Jtsiu6 = (~(Ar1iu6 & Fkfpw6[12]));
assign Ctsiu6 = (~(HRDATA[12] & St1iu6));
assign Kqsiu6 = (Qtsiu6 & Xtsiu6);
assign Xtsiu6 = (Eusiu6 & Lusiu6);
assign Lusiu6 = (~(K7hpw6[12] & Kw1iu6));
assign Eusiu6 = (Susiu6 & Zusiu6);
assign Zusiu6 = (~(Gqgpw6[12] & Xs1iu6));
assign Susiu6 = (~(Trgpw6[12] & Dw1iu6));
assign Qtsiu6 = (Gvsiu6 & Nvsiu6);
assign Gvsiu6 = (Uvsiu6 & Bwsiu6);
assign Bwsiu6 = (~(vis_pc_o[11] & Iv1iu6));
assign Ipsiu6 = (Iwsiu6 & Pwsiu6);
assign Pwsiu6 = (~(Jshpw6[12] & Bo1iu6));
assign Iwsiu6 = (~(Uthpw6[12] & Sf1iu6));
assign Hbphu6 = (~(Wwsiu6 & Dxsiu6));
assign Dxsiu6 = (Kxsiu6 & Po1iu6);
assign Kxsiu6 = (~(Wo1iu6 & Rxsiu6));
assign Rxsiu6 = (~(Yxsiu6 & Fysiu6));
assign Fysiu6 = (Mysiu6 & Tysiu6);
assign Tysiu6 = (Azsiu6 & Hzsiu6);
assign Hzsiu6 = (~(Ar1iu6 & Fkfpw6[13]));
assign Azsiu6 = (Ozsiu6 & Vzsiu6);
assign Vzsiu6 = (~(Togpw6[13] & Vr1iu6));
assign Ozsiu6 = (~(Gtgpw6[13] & Cs1iu6));
assign Mysiu6 = (C0tiu6 & J0tiu6);
assign J0tiu6 = (~(Gqgpw6[13] & Xs1iu6));
assign C0tiu6 = (Q0tiu6 & X0tiu6);
assign X0tiu6 = (~(HRDATA[13] & St1iu6));
assign Q0tiu6 = (~(E1hpw6[13] & Zt1iu6));
assign Yxsiu6 = (E1tiu6 & L1tiu6);
assign L1tiu6 = (S1tiu6 & Z1tiu6);
assign Z1tiu6 = (~(vis_pc_o[12] & Iv1iu6));
assign S1tiu6 = (G2tiu6 & N2tiu6);
assign N2tiu6 = (~(Trgpw6[13] & Dw1iu6));
assign G2tiu6 = (~(K7hpw6[13] & Kw1iu6));
assign E1tiu6 = (U2tiu6 & Yw1iu6);
assign Wwsiu6 = (B3tiu6 & I3tiu6);
assign I3tiu6 = (~(Jshpw6[13] & Bo1iu6));
assign B3tiu6 = (~(Uthpw6[13] & Sf1iu6));
assign Abphu6 = (~(P3tiu6 & W3tiu6));
assign W3tiu6 = (D4tiu6 & Po1iu6);
assign D4tiu6 = (~(Wo1iu6 & K4tiu6));
assign K4tiu6 = (~(R4tiu6 & Y4tiu6));
assign Y4tiu6 = (F5tiu6 & M5tiu6);
assign M5tiu6 = (T5tiu6 & A6tiu6);
assign A6tiu6 = (~(Ar1iu6 & Fkfpw6[14]));
assign T5tiu6 = (H6tiu6 & O6tiu6);
assign O6tiu6 = (~(Togpw6[14] & Vr1iu6));
assign H6tiu6 = (~(Gtgpw6[14] & Cs1iu6));
assign F5tiu6 = (V6tiu6 & C7tiu6);
assign C7tiu6 = (~(Gqgpw6[14] & Xs1iu6));
assign V6tiu6 = (J7tiu6 & Q7tiu6);
assign Q7tiu6 = (~(HRDATA[14] & St1iu6));
assign J7tiu6 = (~(E1hpw6[14] & Zt1iu6));
assign R4tiu6 = (X7tiu6 & E8tiu6);
assign E8tiu6 = (L8tiu6 & S8tiu6);
assign S8tiu6 = (~(vis_pc_o[13] & Iv1iu6));
assign L8tiu6 = (Z8tiu6 & G9tiu6);
assign G9tiu6 = (~(Trgpw6[14] & Dw1iu6));
assign Z8tiu6 = (~(K7hpw6[14] & Kw1iu6));
assign X7tiu6 = (N9tiu6 & Uvsiu6);
assign P3tiu6 = (U9tiu6 & Batiu6);
assign Batiu6 = (~(Jshpw6[14] & Bo1iu6));
assign U9tiu6 = (~(Uthpw6[14] & Sf1iu6));
assign Taphu6 = (~(Iatiu6 & Patiu6));
assign Patiu6 = (Watiu6 & Po1iu6);
assign Watiu6 = (~(Wo1iu6 & Dbtiu6));
assign Dbtiu6 = (~(Kbtiu6 & Rbtiu6));
assign Rbtiu6 = (Ybtiu6 & Fctiu6);
assign Fctiu6 = (Mctiu6 & Tctiu6);
assign Tctiu6 = (~(Ar1iu6 & Fkfpw6[15]));
assign Mctiu6 = (Adtiu6 & Hdtiu6);
assign Hdtiu6 = (~(Togpw6[15] & Vr1iu6));
assign Adtiu6 = (~(Gtgpw6[15] & Cs1iu6));
assign Ybtiu6 = (Odtiu6 & Vdtiu6);
assign Vdtiu6 = (~(Gqgpw6[15] & Xs1iu6));
assign Odtiu6 = (Cetiu6 & Jetiu6);
assign Jetiu6 = (~(HRDATA[15] & St1iu6));
assign Cetiu6 = (~(E1hpw6[15] & Zt1iu6));
assign Kbtiu6 = (Qetiu6 & Xetiu6);
assign Xetiu6 = (Eftiu6 & Lftiu6);
assign Lftiu6 = (~(vis_pc_o[14] & Iv1iu6));
assign Eftiu6 = (Sftiu6 & Zftiu6);
assign Zftiu6 = (~(Trgpw6[15] & Dw1iu6));
assign Sftiu6 = (~(K7hpw6[15] & Kw1iu6));
assign Qetiu6 = (Ggtiu6 & Uvsiu6);
assign Iatiu6 = (Ngtiu6 & Ugtiu6);
assign Ugtiu6 = (~(Jshpw6[15] & Bo1iu6));
assign Ngtiu6 = (~(Uthpw6[15] & Sf1iu6));
assign Maphu6 = (~(Bhtiu6 & Ihtiu6));
assign Ihtiu6 = (Phtiu6 & Whtiu6);
assign Whtiu6 = (~(Wo1iu6 & Ditiu6));
assign Ditiu6 = (~(Kitiu6 & Ritiu6));
assign Ritiu6 = (Yitiu6 & Fjtiu6);
assign Fjtiu6 = (Mjtiu6 & Tjtiu6);
assign Tjtiu6 = (~(Ar1iu6 & Fkfpw6[16]));
assign Mjtiu6 = (Aktiu6 & Hktiu6);
assign Hktiu6 = (~(Togpw6[16] & Vr1iu6));
assign Aktiu6 = (~(Gtgpw6[16] & Cs1iu6));
assign Yitiu6 = (Oktiu6 & Vktiu6);
assign Vktiu6 = (~(Gqgpw6[16] & Xs1iu6));
assign Oktiu6 = (Cltiu6 & Jltiu6);
assign Jltiu6 = (~(HRDATA[16] & St1iu6));
assign Cltiu6 = (~(E1hpw6[16] & Zt1iu6));
assign Kitiu6 = (Qltiu6 & Xltiu6);
assign Xltiu6 = (Emtiu6 & Lmtiu6);
assign Lmtiu6 = (~(vis_pc_o[15] & Iv1iu6));
assign Emtiu6 = (Smtiu6 & Zmtiu6);
assign Zmtiu6 = (~(Trgpw6[16] & Dw1iu6));
assign Smtiu6 = (~(K7hpw6[16] & Kw1iu6));
assign Qltiu6 = (Gntiu6 & Nntiu6);
assign Phtiu6 = (~(Jshpw6[16] & Bo1iu6));
assign Bhtiu6 = (Untiu6 & Botiu6);
assign Botiu6 = (~(Uthpw6[16] & Sf1iu6));
assign Faphu6 = (~(Iotiu6 & Potiu6));
assign Potiu6 = (Wotiu6 & Dptiu6);
assign Dptiu6 = (~(Wo1iu6 & Kptiu6));
assign Kptiu6 = (~(Rptiu6 & Yptiu6));
assign Yptiu6 = (Fqtiu6 & Mqtiu6);
assign Mqtiu6 = (Tqtiu6 & Artiu6);
assign Artiu6 = (~(Ar1iu6 & Fkfpw6[17]));
assign Tqtiu6 = (Hrtiu6 & Ortiu6);
assign Ortiu6 = (~(Togpw6[17] & Vr1iu6));
assign Hrtiu6 = (~(Gtgpw6[17] & Cs1iu6));
assign Fqtiu6 = (Vrtiu6 & Cstiu6);
assign Cstiu6 = (~(Gqgpw6[17] & Xs1iu6));
assign Vrtiu6 = (Jstiu6 & Qstiu6);
assign Qstiu6 = (~(HRDATA[17] & St1iu6));
assign Jstiu6 = (~(E1hpw6[17] & Zt1iu6));
assign Rptiu6 = (Xstiu6 & Ettiu6);
assign Ettiu6 = (Lttiu6 & Sttiu6);
assign Sttiu6 = (~(vis_pc_o[16] & Iv1iu6));
assign Lttiu6 = (Zttiu6 & Gutiu6);
assign Gutiu6 = (~(Trgpw6[17] & Dw1iu6));
assign Zttiu6 = (~(K7hpw6[17] & Kw1iu6));
assign Xstiu6 = (Nutiu6 & Nntiu6);
assign Nntiu6 = (Reqiu6 & Uutiu6);
assign Uutiu6 = (~(HALTED & Bvtiu6));
assign Wotiu6 = (~(Jshpw6[17] & Bo1iu6));
assign Iotiu6 = (Untiu6 & Ivtiu6);
assign Ivtiu6 = (~(Uthpw6[17] & Sf1iu6));
assign Y9phu6 = (~(Pvtiu6 & Wvtiu6));
assign Wvtiu6 = (Dwtiu6 & Kwtiu6);
assign Kwtiu6 = (~(Wo1iu6 & Rwtiu6));
assign Rwtiu6 = (~(Ywtiu6 & Fxtiu6));
assign Fxtiu6 = (Mxtiu6 & Txtiu6);
assign Txtiu6 = (Aytiu6 & Hytiu6);
assign Hytiu6 = (Duhiu6 | Qa5iu6);
assign Aytiu6 = (Oytiu6 & Reqiu6);
assign Oytiu6 = (~(Togpw6[18] & Vr1iu6));
assign Mxtiu6 = (Vytiu6 & Cztiu6);
assign Cztiu6 = (~(HRDATA[18] & St1iu6));
assign Vytiu6 = (Jztiu6 & Qztiu6);
assign Qztiu6 = (~(Gtgpw6[18] & Cs1iu6));
assign Jztiu6 = (~(Ar1iu6 & Fkfpw6[18]));
assign Ywtiu6 = (Xztiu6 & E0uiu6);
assign E0uiu6 = (L0uiu6 & S0uiu6);
assign S0uiu6 = (~(Trgpw6[18] & Dw1iu6));
assign L0uiu6 = (Z0uiu6 & G1uiu6);
assign G1uiu6 = (~(E1hpw6[18] & Zt1iu6));
assign Z0uiu6 = (~(Gqgpw6[18] & Xs1iu6));
assign Xztiu6 = (N1uiu6 & U1uiu6);
assign N1uiu6 = (B2uiu6 & I2uiu6);
assign I2uiu6 = (~(K7hpw6[18] & Kw1iu6));
assign B2uiu6 = (~(vis_pc_o[17] & Iv1iu6));
assign Dwtiu6 = (~(Jshpw6[18] & Bo1iu6));
assign Pvtiu6 = (Untiu6 & P2uiu6);
assign P2uiu6 = (~(Uthpw6[18] & Sf1iu6));
assign R9phu6 = (~(W2uiu6 & D3uiu6));
assign D3uiu6 = (K3uiu6 & Po1iu6);
assign K3uiu6 = (~(Wo1iu6 & R3uiu6));
assign R3uiu6 = (~(Y3uiu6 & F4uiu6));
assign F4uiu6 = (M4uiu6 & T4uiu6);
assign T4uiu6 = (A5uiu6 & H5uiu6);
assign H5uiu6 = (Duhiu6 | Dp8iu6);
assign A5uiu6 = (O5uiu6 & Reqiu6);
assign O5uiu6 = (~(Togpw6[19] & Vr1iu6));
assign M4uiu6 = (V5uiu6 & C6uiu6);
assign C6uiu6 = (~(HRDATA[19] & St1iu6));
assign V5uiu6 = (J6uiu6 & Q6uiu6);
assign Q6uiu6 = (~(Gtgpw6[19] & Cs1iu6));
assign J6uiu6 = (~(Ar1iu6 & Fkfpw6[19]));
assign Y3uiu6 = (X6uiu6 & E7uiu6);
assign E7uiu6 = (L7uiu6 & S7uiu6);
assign S7uiu6 = (~(Trgpw6[19] & Dw1iu6));
assign L7uiu6 = (Z7uiu6 & G8uiu6);
assign G8uiu6 = (~(E1hpw6[19] & Zt1iu6));
assign Z7uiu6 = (~(Gqgpw6[19] & Xs1iu6));
assign X6uiu6 = (N8uiu6 & U8uiu6);
assign N8uiu6 = (B9uiu6 & I9uiu6);
assign I9uiu6 = (~(K7hpw6[19] & Kw1iu6));
assign B9uiu6 = (~(vis_pc_o[18] & Iv1iu6));
assign W2uiu6 = (P9uiu6 & W9uiu6);
assign W9uiu6 = (~(Jshpw6[19] & Bo1iu6));
assign P9uiu6 = (~(Uthpw6[19] & Sf1iu6));
assign K9phu6 = (~(Dauiu6 & Kauiu6));
assign Kauiu6 = (Rauiu6 & V1riu6);
assign Rauiu6 = (~(Wo1iu6 & Yauiu6));
assign Yauiu6 = (~(Fbuiu6 & Mbuiu6));
assign Mbuiu6 = (Tbuiu6 & Acuiu6);
assign Acuiu6 = (Hcuiu6 & Ocuiu6);
assign Ocuiu6 = (~(Ar1iu6 & Fkfpw6[20]));
assign Hcuiu6 = (Vcuiu6 & Cduiu6);
assign Cduiu6 = (~(Togpw6[20] & Vr1iu6));
assign Vcuiu6 = (~(Gtgpw6[20] & Cs1iu6));
assign Tbuiu6 = (Jduiu6 & Qduiu6);
assign Qduiu6 = (~(Gqgpw6[20] & Xs1iu6));
assign Jduiu6 = (Xduiu6 & Eeuiu6);
assign Eeuiu6 = (~(HRDATA[20] & St1iu6));
assign Xduiu6 = (~(E1hpw6[20] & Zt1iu6));
assign Fbuiu6 = (Leuiu6 & Seuiu6);
assign Seuiu6 = (Zeuiu6 & Gfuiu6);
assign Gfuiu6 = (~(vis_pc_o[19] & Iv1iu6));
assign Zeuiu6 = (Nfuiu6 & Ufuiu6);
assign Ufuiu6 = (~(Trgpw6[20] & Dw1iu6));
assign Nfuiu6 = (~(K7hpw6[20] & Kw1iu6));
assign Leuiu6 = (Bguiu6 & Yw1iu6);
assign Dauiu6 = (Iguiu6 & Pguiu6);
assign Pguiu6 = (~(Jshpw6[20] & Bo1iu6));
assign Iguiu6 = (~(Uthpw6[20] & Sf1iu6));
assign D9phu6 = (~(Wguiu6 & Dhuiu6));
assign Dhuiu6 = (Khuiu6 & V1riu6);
assign Khuiu6 = (~(Wo1iu6 & Rhuiu6));
assign Rhuiu6 = (~(Yhuiu6 & Fiuiu6));
assign Fiuiu6 = (Miuiu6 & Tiuiu6);
assign Tiuiu6 = (Ajuiu6 & Hjuiu6);
assign Hjuiu6 = (~(Ar1iu6 & Fkfpw6[21]));
assign Ajuiu6 = (Ojuiu6 & Vjuiu6);
assign Vjuiu6 = (~(Togpw6[21] & Vr1iu6));
assign Ojuiu6 = (~(Gtgpw6[21] & Cs1iu6));
assign Miuiu6 = (Ckuiu6 & Jkuiu6);
assign Jkuiu6 = (~(Gqgpw6[21] & Xs1iu6));
assign Ckuiu6 = (Qkuiu6 & Xkuiu6);
assign Xkuiu6 = (~(HRDATA[21] & St1iu6));
assign Qkuiu6 = (~(E1hpw6[21] & Zt1iu6));
assign Yhuiu6 = (Eluiu6 & Lluiu6);
assign Lluiu6 = (Sluiu6 & Zluiu6);
assign Zluiu6 = (~(vis_pc_o[20] & Iv1iu6));
assign Sluiu6 = (Gmuiu6 & Nmuiu6);
assign Nmuiu6 = (~(Trgpw6[21] & Dw1iu6));
assign Gmuiu6 = (~(K7hpw6[21] & Kw1iu6));
assign Eluiu6 = (Umuiu6 & Yw1iu6);
assign Wguiu6 = (Bnuiu6 & Inuiu6);
assign Inuiu6 = (~(Jshpw6[21] & Bo1iu6));
assign Bnuiu6 = (~(Uthpw6[21] & Sf1iu6));
assign W8phu6 = (~(Pnuiu6 & Wnuiu6));
assign Wnuiu6 = (Douiu6 & V1riu6);
assign Douiu6 = (~(Wo1iu6 & Kouiu6));
assign Kouiu6 = (~(Rouiu6 & Youiu6));
assign Youiu6 = (Fpuiu6 & Mpuiu6);
assign Mpuiu6 = (Tpuiu6 & Aquiu6);
assign Aquiu6 = (~(Ar1iu6 & Fkfpw6[22]));
assign Tpuiu6 = (Hquiu6 & Oquiu6);
assign Oquiu6 = (~(Togpw6[22] & Vr1iu6));
assign Hquiu6 = (~(Gtgpw6[22] & Cs1iu6));
assign Fpuiu6 = (Vquiu6 & Cruiu6);
assign Cruiu6 = (~(Gqgpw6[22] & Xs1iu6));
assign Vquiu6 = (Jruiu6 & Qruiu6);
assign Qruiu6 = (~(HRDATA[22] & St1iu6));
assign Jruiu6 = (~(E1hpw6[22] & Zt1iu6));
assign Rouiu6 = (Xruiu6 & Esuiu6);
assign Esuiu6 = (Lsuiu6 & Ssuiu6);
assign Ssuiu6 = (~(vis_pc_o[21] & Iv1iu6));
assign Lsuiu6 = (Zsuiu6 & Gtuiu6);
assign Gtuiu6 = (~(Trgpw6[22] & Dw1iu6));
assign Zsuiu6 = (~(K7hpw6[22] & Kw1iu6));
assign Xruiu6 = (Ntuiu6 & Yw1iu6);
assign Pnuiu6 = (Utuiu6 & Buuiu6);
assign Buuiu6 = (~(Jshpw6[22] & Bo1iu6));
assign Utuiu6 = (~(Uthpw6[22] & Sf1iu6));
assign P8phu6 = (~(Iuuiu6 & Puuiu6));
assign Puuiu6 = (~(Uthpw6[23] & Sf1iu6));
assign Iuuiu6 = (Wuuiu6 & Dvuiu6);
assign Dvuiu6 = (~(Wo1iu6 & Kvuiu6));
assign Kvuiu6 = (~(Rvuiu6 & Yvuiu6));
assign Yvuiu6 = (Fwuiu6 & Mwuiu6);
assign Mwuiu6 = (Twuiu6 & Axuiu6);
assign Axuiu6 = (~(Ar1iu6 & Fkfpw6[23]));
assign Twuiu6 = (Hxuiu6 & Oxuiu6);
assign Oxuiu6 = (~(Togpw6[23] & Vr1iu6));
assign Hxuiu6 = (~(Gtgpw6[23] & Cs1iu6));
assign Fwuiu6 = (Vxuiu6 & Cyuiu6);
assign Cyuiu6 = (~(Gqgpw6[23] & Xs1iu6));
assign Vxuiu6 = (Jyuiu6 & Qyuiu6);
assign Qyuiu6 = (~(HRDATA[23] & St1iu6));
assign Jyuiu6 = (~(E1hpw6[23] & Zt1iu6));
assign Rvuiu6 = (Xyuiu6 & Ezuiu6);
assign Ezuiu6 = (Lzuiu6 & Szuiu6);
assign Szuiu6 = (~(vis_pc_o[22] & Iv1iu6));
assign Lzuiu6 = (Zzuiu6 & G0viu6);
assign G0viu6 = (~(Trgpw6[23] & Dw1iu6));
assign Zzuiu6 = (~(K7hpw6[23] & Kw1iu6));
assign Xyuiu6 = (N0viu6 & Yw1iu6);
assign Wuuiu6 = (~(Jshpw6[23] & Bo1iu6));
assign I8phu6 = (~(U0viu6 & B1viu6));
assign B1viu6 = (I1viu6 & Bcriu6);
assign I1viu6 = (~(Wo1iu6 & P1viu6));
assign P1viu6 = (~(W1viu6 & D2viu6));
assign D2viu6 = (K2viu6 & R2viu6);
assign R2viu6 = (Y2viu6 & F3viu6);
assign F3viu6 = (M3viu6 & T3viu6);
assign T3viu6 = (~(Vxmhu6 & Eg7iu6));
assign M3viu6 = (~(Yc7iu6 & E5hhu6));
assign Y2viu6 = (A4viu6 & H4viu6);
assign H4viu6 = (~(Togpw6[24] & Vr1iu6));
assign A4viu6 = (~(R6hhu6 & Bvtiu6));
assign K2viu6 = (O4viu6 & V4viu6);
assign V4viu6 = (C5viu6 & J5viu6);
assign J5viu6 = (~(Hwmhu6 & Ws4iu6));
assign C5viu6 = (~(Gtgpw6[24] & Cs1iu6));
assign O4viu6 = (Q5viu6 & X5viu6);
assign X5viu6 = (~(Ar1iu6 & Fkfpw6[24]));
assign Q5viu6 = (~(HRDATA[24] & St1iu6));
assign W1viu6 = (E6viu6 & L6viu6);
assign L6viu6 = (S6viu6 & Z6viu6);
assign Z6viu6 = (G7viu6 & N7viu6);
assign N7viu6 = (~(E1hpw6[24] & Zt1iu6));
assign G7viu6 = (~(Gqgpw6[24] & Xs1iu6));
assign S6viu6 = (U7viu6 & B8viu6);
assign B8viu6 = (~(Trgpw6[24] & Dw1iu6));
assign U7viu6 = (~(K7hpw6[24] & Kw1iu6));
assign E6viu6 = (I8viu6 & P8viu6);
assign I8viu6 = (Yw1iu6 & W8viu6);
assign W8viu6 = (~(vis_pc_o[23] & Iv1iu6));
assign U0viu6 = (D9viu6 & K9viu6);
assign K9viu6 = (~(Jshpw6[24] & Bo1iu6));
assign D9viu6 = (~(Uthpw6[24] & Sf1iu6));
assign B8phu6 = (~(R9viu6 & Y9viu6));
assign Y9viu6 = (Faviu6 & Bcriu6);
assign Bcriu6 = (!Qwpiu6);
assign Faviu6 = (~(Wo1iu6 & Maviu6));
assign Maviu6 = (~(Taviu6 & Abviu6));
assign Abviu6 = (Hbviu6 & Obviu6);
assign Obviu6 = (Vbviu6 & Ccviu6);
assign Ccviu6 = (~(Gtgpw6[25] & Cs1iu6));
assign Vbviu6 = (Jcviu6 & Qcviu6);
assign Qcviu6 = (~(Togpw6[25] & Vr1iu6));
assign Jcviu6 = (~(D8hhu6 & Bvtiu6));
assign Hbviu6 = (Xcviu6 & Edviu6);
assign Edviu6 = (~(E1hpw6[25] & Zt1iu6));
assign Xcviu6 = (Ldviu6 & Sdviu6);
assign Sdviu6 = (~(Ar1iu6 & Fkfpw6[25]));
assign Ldviu6 = (~(HRDATA[25] & St1iu6));
assign Taviu6 = (Zdviu6 & Geviu6);
assign Geviu6 = (Neviu6 & Ueviu6);
assign Ueviu6 = (~(K7hpw6[25] & Kw1iu6));
assign Neviu6 = (Bfviu6 & Ifviu6);
assign Ifviu6 = (~(Gqgpw6[25] & Xs1iu6));
assign Bfviu6 = (~(Trgpw6[25] & Dw1iu6));
assign Zdviu6 = (Pfviu6 & Wfviu6);
assign Pfviu6 = (Yw1iu6 & Dgviu6);
assign Dgviu6 = (~(vis_pc_o[24] & Iv1iu6));
assign R9viu6 = (Kgviu6 & Rgviu6);
assign Rgviu6 = (~(Jshpw6[25] & Bo1iu6));
assign Kgviu6 = (~(Uthpw6[25] & Sf1iu6));
assign U7phu6 = (~(Ygviu6 & Fhviu6));
assign Fhviu6 = (Mhviu6 & V1riu6);
assign Mhviu6 = (~(Wo1iu6 & Thviu6));
assign Thviu6 = (~(Aiviu6 & Hiviu6));
assign Hiviu6 = (Oiviu6 & Viviu6);
assign Viviu6 = (Cjviu6 & Jjviu6);
assign Jjviu6 = (~(Ar1iu6 & Fkfpw6[26]));
assign Cjviu6 = (Qjviu6 & Xjviu6);
assign Xjviu6 = (~(Togpw6[26] & Vr1iu6));
assign Qjviu6 = (~(Gtgpw6[26] & Cs1iu6));
assign Oiviu6 = (Ekviu6 & Lkviu6);
assign Lkviu6 = (~(Gqgpw6[26] & Xs1iu6));
assign Ekviu6 = (Skviu6 & Zkviu6);
assign Zkviu6 = (~(HRDATA[26] & St1iu6));
assign Skviu6 = (~(E1hpw6[26] & Zt1iu6));
assign Aiviu6 = (Glviu6 & Nlviu6);
assign Nlviu6 = (Ulviu6 & Bmviu6);
assign Bmviu6 = (~(vis_pc_o[25] & Iv1iu6));
assign Ulviu6 = (Imviu6 & Pmviu6);
assign Pmviu6 = (~(Trgpw6[26] & Dw1iu6));
assign Imviu6 = (~(K7hpw6[26] & Kw1iu6));
assign Glviu6 = (Wmviu6 & Yw1iu6);
assign Ygviu6 = (Dnviu6 & Knviu6);
assign Knviu6 = (~(Jshpw6[26] & Bo1iu6));
assign Dnviu6 = (~(Uthpw6[26] & Sf1iu6));
assign N7phu6 = (~(Rnviu6 & Ynviu6));
assign Ynviu6 = (~(Uthpw6[27] & Sf1iu6));
assign Rnviu6 = (Foviu6 & Moviu6);
assign Moviu6 = (~(Wo1iu6 & Toviu6));
assign Toviu6 = (~(Apviu6 & Hpviu6));
assign Hpviu6 = (Opviu6 & Vpviu6);
assign Vpviu6 = (Cqviu6 & Jqviu6);
assign Jqviu6 = (~(Ar1iu6 & Fkfpw6[27]));
assign Cqviu6 = (Qqviu6 & Xqviu6);
assign Xqviu6 = (~(Togpw6[27] & Vr1iu6));
assign Qqviu6 = (~(Gtgpw6[27] & Cs1iu6));
assign Opviu6 = (Erviu6 & Lrviu6);
assign Lrviu6 = (~(Gqgpw6[27] & Xs1iu6));
assign Erviu6 = (Srviu6 & Zrviu6);
assign Zrviu6 = (~(HRDATA[27] & St1iu6));
assign Srviu6 = (~(E1hpw6[27] & Zt1iu6));
assign Apviu6 = (Gsviu6 & Nsviu6);
assign Nsviu6 = (Usviu6 & Btviu6);
assign Btviu6 = (~(vis_pc_o[26] & Iv1iu6));
assign Usviu6 = (Itviu6 & Ptviu6);
assign Ptviu6 = (~(Trgpw6[27] & Dw1iu6));
assign Itviu6 = (~(K7hpw6[27] & Kw1iu6));
assign Gsviu6 = (Wtviu6 & Yw1iu6);
assign Foviu6 = (~(Jshpw6[27] & Bo1iu6));
assign G7phu6 = (~(Duviu6 & Kuviu6));
assign Kuviu6 = (Ruviu6 & Yuviu6);
assign Yuviu6 = (~(Wo1iu6 & Fvviu6));
assign Fvviu6 = (~(Mvviu6 & Tvviu6));
assign Tvviu6 = (Awviu6 & Hwviu6);
assign Hwviu6 = (Owviu6 & Vwviu6);
assign Vwviu6 = (~(Ar1iu6 & Fkfpw6[28]));
assign Owviu6 = (Cxviu6 & Jxviu6);
assign Jxviu6 = (~(Togpw6[28] & Vr1iu6));
assign Cxviu6 = (~(Gtgpw6[28] & Cs1iu6));
assign Awviu6 = (Qxviu6 & Xxviu6);
assign Xxviu6 = (~(Gqgpw6[28] & Xs1iu6));
assign Qxviu6 = (Eyviu6 & Lyviu6);
assign Lyviu6 = (~(HRDATA[28] & St1iu6));
assign Eyviu6 = (~(E1hpw6[28] & Zt1iu6));
assign Mvviu6 = (Syviu6 & Zyviu6);
assign Zyviu6 = (Gzviu6 & Nzviu6);
assign Nzviu6 = (~(Iv1iu6 & vis_pc_o[27]));
assign Gzviu6 = (Uzviu6 & B0wiu6);
assign B0wiu6 = (~(Trgpw6[28] & Dw1iu6));
assign Uzviu6 = (~(K7hpw6[28] & Kw1iu6));
assign Syviu6 = (I0wiu6 & Yw1iu6);
assign Ruviu6 = (~(Jshpw6[28] & Bo1iu6));
assign Duviu6 = (P0wiu6 & W0wiu6);
assign W0wiu6 = (~(ECOREVNUM[20] & Tx1iu6));
assign P0wiu6 = (~(Uthpw6[28] & Sf1iu6));
assign Z6phu6 = (~(D1wiu6 & K1wiu6));
assign K1wiu6 = (R1wiu6 & Y1wiu6);
assign Y1wiu6 = (~(Jshpw6[29] & Bo1iu6));
assign R1wiu6 = (F2wiu6 & Po1iu6);
assign F2wiu6 = (~(Wo1iu6 & M2wiu6));
assign M2wiu6 = (~(T2wiu6 & A3wiu6));
assign A3wiu6 = (H3wiu6 & O3wiu6);
assign O3wiu6 = (V3wiu6 & C4wiu6);
assign C4wiu6 = (~(J4wiu6 & C3qiu6));
assign J4wiu6 = (Q4wiu6 & X4wiu6);
assign V3wiu6 = (~(Ar1iu6 & Fkfpw6[29]));
assign H3wiu6 = (E5wiu6 & L5wiu6);
assign L5wiu6 = (~(HRDATA[29] & St1iu6));
assign E5wiu6 = (~(E1hpw6[29] & Zt1iu6));
assign T2wiu6 = (S5wiu6 & Z5wiu6);
assign Z5wiu6 = (G6wiu6 & N6wiu6);
assign N6wiu6 = (~(K7hpw6[29] & Kw1iu6));
assign G6wiu6 = (~(Iv1iu6 & vis_pc_o[28]));
assign S5wiu6 = (U6wiu6 & Yw1iu6);
assign D1wiu6 = (B7wiu6 & I7wiu6);
assign I7wiu6 = (~(ECOREVNUM[21] & Tx1iu6));
assign B7wiu6 = (~(Uthpw6[29] & Sf1iu6));
assign S6phu6 = (~(P7wiu6 & W7wiu6));
assign W7wiu6 = (D8wiu6 & K8wiu6);
assign K8wiu6 = (~(Jshpw6[30] & Bo1iu6));
assign D8wiu6 = (R8wiu6 & Po1iu6);
assign R8wiu6 = (~(Wo1iu6 & Y8wiu6));
assign Y8wiu6 = (~(F9wiu6 & M9wiu6));
assign M9wiu6 = (T9wiu6 & Aawiu6);
assign Aawiu6 = (Hawiu6 & Oawiu6);
assign Oawiu6 = (~(Ar1iu6 & Fkfpw6[30]));
assign Hawiu6 = (Vawiu6 & Cbwiu6);
assign Cbwiu6 = (~(Ligpw6[27] & Vr1iu6));
assign Vawiu6 = (~(Engpw6[27] & Cs1iu6));
assign T9wiu6 = (Jbwiu6 & Qbwiu6);
assign Qbwiu6 = (~(Akgpw6[27] & Xs1iu6));
assign Jbwiu6 = (Xbwiu6 & Ecwiu6);
assign Ecwiu6 = (~(HRDATA[30] & St1iu6));
assign Xbwiu6 = (~(E1hpw6[30] & Zt1iu6));
assign F9wiu6 = (Lcwiu6 & Scwiu6);
assign Scwiu6 = (Zcwiu6 & Gdwiu6);
assign Gdwiu6 = (~(Iv1iu6 & vis_pc_o[29]));
assign Zcwiu6 = (Ndwiu6 & Udwiu6);
assign Udwiu6 = (~(Plgpw6[27] & Dw1iu6));
assign Ndwiu6 = (~(K7hpw6[30] & Kw1iu6));
assign Lcwiu6 = (Bewiu6 & Yw1iu6);
assign P7wiu6 = (Iewiu6 & Pewiu6);
assign Pewiu6 = (~(ECOREVNUM[22] & Tx1iu6));
assign Iewiu6 = (~(Uthpw6[30] & Sf1iu6));
assign L6phu6 = (~(Wewiu6 & Dfwiu6));
assign Dfwiu6 = (Kfwiu6 & Rfwiu6);
assign Rfwiu6 = (~(Qwpiu6 & Aphpw6[1]));
assign Qwpiu6 = (~(Yfwiu6 | Vo4iu6));
assign Kfwiu6 = (Fgwiu6 & Mgwiu6);
assign Mgwiu6 = (~(Tnhpw6[0] & Bo1iu6));
assign Bo1iu6 = (Tgwiu6 & Vo4iu6);
assign Tgwiu6 = (!Yfwiu6);
assign Yfwiu6 = (~(Ahwiu6 & Hhwiu6));
assign Hhwiu6 = (~(Wu9iu6 | Ho4iu6));
assign Ahwiu6 = (~(Ohwiu6 | Sf1iu6));
assign Fgwiu6 = (~(Wo1iu6 & Vhwiu6));
assign Vhwiu6 = (~(Ciwiu6 & Jiwiu6));
assign Jiwiu6 = (Qiwiu6 & Xiwiu6);
assign Xiwiu6 = (Ejwiu6 & Ljwiu6);
assign Ljwiu6 = (Sjwiu6 & Zjwiu6);
assign Zjwiu6 = (~(Gkwiu6 & A2qiu6));
assign Gkwiu6 = (Nkwiu6 & Ukwiu6);
assign Sjwiu6 = (~(Q3qiu6 | U4riu6));
assign U4riu6 = (Ffqiu6 & C3qiu6);
assign Q3qiu6 = (Blwiu6 & X8hpw6[1]);
assign Blwiu6 = (Nkwiu6 & Ilwiu6);
assign Ejwiu6 = (Plwiu6 & Wlwiu6);
assign Wlwiu6 = (~(G4hpw6[0] & Sg7iu6));
assign Sg7iu6 = (Dmwiu6 & Q4wiu6);
assign Plwiu6 = (Kmwiu6 & Rmwiu6);
assign Rmwiu6 = (~(R2hpw6[0] & Eg7iu6));
assign Eg7iu6 = (Vuciu6 & Nkwiu6);
assign Kmwiu6 = (~(Dhgpw6[0] & Fgpiu6));
assign Fgpiu6 = (Ymwiu6 & Fnwiu6);
assign Ymwiu6 = (Mnwiu6 & Ilwiu6);
assign Qiwiu6 = (Tnwiu6 & Aowiu6);
assign Aowiu6 = (Howiu6 & Oowiu6);
assign Oowiu6 = (~(Kohhu6 & Ve7iu6));
assign Ve7iu6 = (Vowiu6 & Cpwiu6);
assign Howiu6 = (Jpwiu6 & Qpwiu6);
assign Qpwiu6 = (~(Yc7iu6 & H2hhu6));
assign Yc7iu6 = (Xpwiu6 & Dzqiu6);
assign Xpwiu6 = (Q4wiu6 & Cvciu6);
assign Jpwiu6 = (~(Aygpw6[0] & Jf7iu6));
assign Jf7iu6 = (Dmwiu6 & Mnwiu6);
assign Dmwiu6 = (Eqwiu6 & C3qiu6);
assign Tnwiu6 = (Lqwiu6 & Sqwiu6);
assign Sqwiu6 = (~(Lwgpw6[0] & Ws4iu6));
assign Ws4iu6 = (~(Zqwiu6 | Mfqiu6));
assign Lqwiu6 = (Grwiu6 & Nrwiu6);
assign Nrwiu6 = (~(Qhhhu6 & Vr1iu6));
assign Vr1iu6 = (Vuciu6 & Urwiu6);
assign Grwiu6 = (Duhiu6 | Zwciu6);
assign Duhiu6 = (!Bvtiu6);
assign Bvtiu6 = (Fnwiu6 & Vuciu6);
assign Fnwiu6 = (Bswiu6 & Dr6iu6);
assign Ciwiu6 = (Iswiu6 & Pswiu6);
assign Pswiu6 = (Wswiu6 & Dtwiu6);
assign Dtwiu6 = (Ktwiu6 & Rtwiu6);
assign Rtwiu6 = (~(HRDATA[0] & St1iu6));
assign St1iu6 = (Ytwiu6 & Ur4iu6);
assign Ur4iu6 = (Fuwiu6 & Q4wiu6);
assign Fuwiu6 = (Cvciu6 & Ukwiu6);
assign Ktwiu6 = (Muwiu6 & Tuwiu6);
assign Tuwiu6 = (~(Smhhu6 & Cs1iu6));
assign Cs1iu6 = (Cpwiu6 & Avwiu6);
assign Muwiu6 = (~(Ar1iu6 & Fkfpw6[0]));
assign Ar1iu6 = (Rzciu6 & D5eiu6);
assign Wswiu6 = (Hvwiu6 & Ovwiu6);
assign Ovwiu6 = (~(Alhhu6 & Dw1iu6));
assign Dw1iu6 = (Avwiu6 & Urwiu6);
assign Urwiu6 = (Vvwiu6 & X8hpw6[6]);
assign Vvwiu6 = (~(X8hpw6[0] | X8hpw6[5]));
assign Hvwiu6 = (Cwwiu6 & Jwwiu6);
assign Jwwiu6 = (~(Zt1iu6 & Pzgpw6[0]));
assign Zt1iu6 = (Avwiu6 & Nkwiu6);
assign Avwiu6 = (Dzqiu6 & Mnwiu6);
assign Cwwiu6 = (~(Ijhhu6 & Xs1iu6));
assign Xs1iu6 = (Cpwiu6 & Vuciu6);
assign Vuciu6 = (Mnwiu6 & Ukwiu6);
assign Iswiu6 = (Qwwiu6 & Xwwiu6);
assign Xwwiu6 = (~(Exwiu6 | Ylqiu6));
assign Ylqiu6 = (~(Lxwiu6 & Sxwiu6));
assign Sxwiu6 = (~(Zxwiu6 & Ffqiu6));
assign Zxwiu6 = (Ilwiu6 & Dr6iu6);
assign Lxwiu6 = (~(Gywiu6 & A2qiu6));
assign Gywiu6 = (Bswiu6 & Nywiu6);
assign Exwiu6 = (~(Yw1iu6 & Uywiu6));
assign Uywiu6 = (~(Kw1iu6 & V5hpw6[0]));
assign Kw1iu6 = (~(Nwriu6 | Zqwiu6));
assign Nwriu6 = (!Dzqiu6);
assign Yw1iu6 = (Bzwiu6 & Uvsiu6);
assign Uvsiu6 = (Izwiu6 & Reqiu6);
assign Reqiu6 = (~(Iv1iu6 & Pzwiu6));
assign Iv1iu6 = (Wzwiu6 & Vowiu6);
assign Vowiu6 = (Q4wiu6 & Ukwiu6);
assign Wzwiu6 = (X8hpw6[0] & Bswiu6);
assign Izwiu6 = (~(D0xiu6 & K0xiu6));
assign D0xiu6 = (Bqriu6 & Q4wiu6);
assign Bzwiu6 = (R0xiu6 & Hssiu6);
assign Hssiu6 = (~(Y0xiu6 & Mnwiu6));
assign Mnwiu6 = (~(Fl6iu6 | X8hpw6[1]));
assign Y0xiu6 = (Ilwiu6 & K0xiu6);
assign R0xiu6 = (Zqwiu6 | J3qiu6);
assign J3qiu6 = (!Bqriu6);
assign Zqwiu6 = (~(Nkwiu6 & Q4wiu6));
assign Qwwiu6 = (F1xiu6 & M1xiu6);
assign F1xiu6 = (Uwriu6 & Qaqiu6);
assign Qaqiu6 = (Anqiu6 & T1xiu6);
assign T1xiu6 = (~(Ffqiu6 & Nywiu6));
assign Nywiu6 = (!A2xiu6);
assign A2xiu6 = (X8hpw6[0] ? Mfqiu6 : H2xiu6);
assign Mfqiu6 = (!Ukwiu6);
assign Ffqiu6 = (O2xiu6 & X8hpw6[1]);
assign O2xiu6 = (Bswiu6 & Fl6iu6);
assign Anqiu6 = (V2xiu6 & C3xiu6);
assign C3xiu6 = (~(Mmqiu6 & A2qiu6));
assign Mmqiu6 = (Nkwiu6 & Bqriu6);
assign Nkwiu6 = (J3xiu6 & X8hpw6[0]);
assign J3xiu6 = (~(Zh6iu6 | X8hpw6[5]));
assign V2xiu6 = (~(Bswiu6 & Q3xiu6));
assign Q3xiu6 = (~(X3xiu6 & E4xiu6));
assign E4xiu6 = (~(Ryriu6 & Dr6iu6));
assign Ryriu6 = (A2qiu6 & L4xiu6);
assign L4xiu6 = (Ilwiu6 | Ukwiu6);
assign X3xiu6 = (~(A2qiu6 & C3qiu6));
assign C3qiu6 = (Dzqiu6 & X8hpw6[0]);
assign A2qiu6 = (X8hpw6[1] & X8hpw6[4]);
assign Bswiu6 = (~(Zh6iu6 | Wj6iu6));
assign Zh6iu6 = (!X8hpw6[6]);
assign Uwriu6 = (S4xiu6 & Z4xiu6);
assign Z4xiu6 = (~(Fl6iu6 & G5xiu6));
assign G5xiu6 = (N5xiu6 | Iqriu6);
assign Iqriu6 = (Ixriu6 & Vm6iu6);
assign Ixriu6 = (U5xiu6 & X8hpw6[1]);
assign U5xiu6 = (K0xiu6 & X8hpw6[2]);
assign K0xiu6 = (Eqwiu6 & X8hpw6[0]);
assign Eqwiu6 = (~(Wj6iu6 | X8hpw6[6]));
assign Wj6iu6 = (!X8hpw6[5]);
assign N5xiu6 = (Wyqiu6 & Ukwiu6);
assign Ukwiu6 = (Eo6iu6 & Vm6iu6);
assign Wyqiu6 = (B6xiu6 & X8hpw6[1]);
assign B6xiu6 = (X8hpw6[0] & X4wiu6);
assign S4xiu6 = (Svriu6 | H2xiu6);
assign H2xiu6 = (~(Bqriu6 | Dzqiu6));
assign Dzqiu6 = (X8hpw6[3] & Eo6iu6);
assign Eo6iu6 = (!X8hpw6[2]);
assign Bqriu6 = (X8hpw6[3] & X8hpw6[2]);
assign Svriu6 = (~(I6xiu6 & X8hpw6[1]));
assign I6xiu6 = (Cvciu6 & Fl6iu6);
assign Fl6iu6 = (!X8hpw6[4]);
assign Cvciu6 = (X4wiu6 & Dr6iu6);
assign Dr6iu6 = (!X8hpw6[0]);
assign X4wiu6 = (~(X8hpw6[5] | X8hpw6[6]));
assign Wo1iu6 = (P6xiu6 & W6xiu6);
assign P6xiu6 = (D7xiu6 & K7xiu6);
assign K7xiu6 = (~(R7xiu6 & Y7xiu6));
assign Y7xiu6 = (Xp4iu6 | C44iu6);
assign D7xiu6 = (!Sf1iu6);
assign Wewiu6 = (Untiu6 & F8xiu6);
assign F8xiu6 = (~(Uthpw6[0] & Sf1iu6));
assign Untiu6 = (V1riu6 & Po1iu6);
assign Po1iu6 = (~(M8xiu6 & C44iu6));
assign V1riu6 = (!Tx1iu6);
assign Tx1iu6 = (M8xiu6 & Vo4iu6);
assign M8xiu6 = (T8xiu6 & A9xiu6);
assign A9xiu6 = (~(R7xiu6 | W6xiu6));
assign W6xiu6 = (!Ohwiu6);
assign Ohwiu6 = (~(Sq4iu6 & H9xiu6));
assign R7xiu6 = (!Ho4iu6);
assign T8xiu6 = (~(Sf1iu6 | Xp4iu6));
assign Xp4iu6 = (!Wu9iu6);
assign Sf1iu6 = (O9xiu6 | Npzhu6);
assign Npzhu6 = (!Sqhpw6[1]);
assign O9xiu6 = (Sqhpw6[0] ? V9xiu6 : Fszhu6);
assign V9xiu6 = (Wqzhu6 | Pqzhu6);
assign Pqzhu6 = (Caxiu6 & Wu9iu6);
assign Wu9iu6 = (Cjhpw6[1] & Iqzhu6);
assign Caxiu6 = (~(C44iu6 | Eq4iu6));
assign C44iu6 = (!Vo4iu6);
assign Vo4iu6 = (Cjhpw6[0] & Iqzhu6);
assign Fszhu6 = (!Drzhu6);
assign Drzhu6 = (HREADY & Jaxiu6);
assign Jaxiu6 = (~(Qaxiu6 & Xaxiu6));
assign Xaxiu6 = (~(HMASTER & Ebxiu6));
assign J5phu6 = (Fk7iu6 & Lbxiu6);
assign Lbxiu6 = (~(Sbxiu6 & Zbxiu6));
assign Zbxiu6 = (~(Xudpw6 & IRQ[0]));
assign Sbxiu6 = (Gcxiu6 & Yj7iu6);
assign Yj7iu6 = (~(Kwfiu6 & HWDATA[0]));
assign Gcxiu6 = (~(Odgpw6[0] & Ncxiu6));
assign Ncxiu6 = (~(K66iu6 & HWDATA[0]));
assign Fk7iu6 = (Sb5iu6 | Ucxiu6);
assign C5phu6 = (Dogiu6 & Bdxiu6);
assign Bdxiu6 = (~(Idxiu6 & Pdxiu6));
assign Pdxiu6 = (~(Fsdpw6 & IRQ[1]));
assign Idxiu6 = (Wdxiu6 & Wngiu6);
assign Wngiu6 = (~(Kwfiu6 & I4eiu6));
assign Wdxiu6 = (~(Odgpw6[1] & Dexiu6));
assign Dexiu6 = (~(K66iu6 & I4eiu6));
assign I4eiu6 = (Npdhu6 & HWDATA[1]);
assign Dogiu6 = (Sb5iu6 | Kexiu6);
assign Kexiu6 = (!Yogiu6);
assign V4phu6 = (Zlgiu6 & Rexiu6);
assign Rexiu6 = (~(Yexiu6 & Ffxiu6));
assign Ffxiu6 = (~(Eodpw6 & IRQ[2]));
assign Yexiu6 = (Mfxiu6 & Slgiu6);
assign Slgiu6 = (~(G3eiu6 & Kwfiu6));
assign Mfxiu6 = (~(Odgpw6[2] & Tfxiu6));
assign Tfxiu6 = (~(G3eiu6 & K66iu6));
assign Zlgiu6 = (Sb5iu6 | Agxiu6);
assign O4phu6 = (Xefiu6 & Hgxiu6);
assign Hgxiu6 = (~(Ogxiu6 & Vgxiu6));
assign Vgxiu6 = (~(Jndpw6 & IRQ[3]));
assign Ogxiu6 = (Chxiu6 & Qefiu6);
assign Qefiu6 = (~(Kwfiu6 & HWDATA[3]));
assign Chxiu6 = (~(Odgpw6[3] & Jhxiu6));
assign Jhxiu6 = (~(K66iu6 & HWDATA[3]));
assign Xefiu6 = (Sb5iu6 | Qhxiu6);
assign H4phu6 = (Tcfiu6 & Xhxiu6);
assign Xhxiu6 = (~(Eixiu6 & Lixiu6));
assign Lixiu6 = (~(Qndpw6 & IRQ[4]));
assign Eixiu6 = (Sixiu6 & Mcfiu6);
assign Mcfiu6 = (~(Kwfiu6 & HWDATA[4]));
assign Sixiu6 = (~(Odgpw6[4] & Zixiu6));
assign Zixiu6 = (~(K66iu6 & HWDATA[4]));
assign Tcfiu6 = (Sb5iu6 | Gjxiu6);
assign Gjxiu6 = (!Odfiu6);
assign A4phu6 = (Pafiu6 & Njxiu6);
assign Njxiu6 = (~(Ujxiu6 & Bkxiu6));
assign Bkxiu6 = (~(Gpdpw6 & IRQ[5]));
assign Ujxiu6 = (Ikxiu6 & Iafiu6);
assign Iafiu6 = (~(Kwfiu6 & HWDATA[5]));
assign Ikxiu6 = (~(Odgpw6[5] & Pkxiu6));
assign Pkxiu6 = (~(K66iu6 & HWDATA[5]));
assign Pafiu6 = (Sb5iu6 | Wkxiu6);
assign T3phu6 = (L8fiu6 & Dlxiu6);
assign Dlxiu6 = (~(Klxiu6 & Rlxiu6));
assign Rlxiu6 = (~(Lodpw6 & IRQ[6]));
assign Klxiu6 = (Ylxiu6 & E8fiu6);
assign E8fiu6 = (~(Kwfiu6 & HWDATA[6]));
assign Ylxiu6 = (~(Odgpw6[6] & Fmxiu6));
assign Fmxiu6 = (~(K66iu6 & HWDATA[6]));
assign L8fiu6 = (Sb5iu6 | Mmxiu6);
assign M3phu6 = (H6fiu6 & Tmxiu6);
assign Tmxiu6 = (~(Anxiu6 & Hnxiu6));
assign Hnxiu6 = (~(Zodpw6 & IRQ[7]));
assign Anxiu6 = (Onxiu6 & A6fiu6);
assign A6fiu6 = (~(Kwfiu6 & HWDATA[7]));
assign Onxiu6 = (~(Odgpw6[7] & Vnxiu6));
assign Vnxiu6 = (~(K66iu6 & HWDATA[7]));
assign H6fiu6 = (Sb5iu6 | Coxiu6);
assign F3phu6 = (Mbgiu6 & Joxiu6);
assign Joxiu6 = (~(Qoxiu6 & Xoxiu6));
assign Xoxiu6 = (~(Judpw6 & IRQ[10]));
assign Qoxiu6 = (Epxiu6 & Fbgiu6);
assign Fbgiu6 = (~(Kwfiu6 & HWDATA[10]));
assign Epxiu6 = (~(Odgpw6[10] & Lpxiu6));
assign Lpxiu6 = (~(K66iu6 & HWDATA[10]));
assign Mbgiu6 = (Sb5iu6 | Spxiu6);
assign Y2phu6 = (I9giu6 & Zpxiu6);
assign Zpxiu6 = (~(Gqxiu6 & Nqxiu6));
assign Nqxiu6 = (~(Cudpw6 & IRQ[11]));
assign Gqxiu6 = (Uqxiu6 & B9giu6);
assign B9giu6 = (~(Kwfiu6 & HWDATA[11]));
assign Uqxiu6 = (~(Odgpw6[11] & Brxiu6));
assign Brxiu6 = (~(K66iu6 & HWDATA[11]));
assign I9giu6 = (Sb5iu6 | Irxiu6);
assign R2phu6 = (E7giu6 & Prxiu6);
assign Prxiu6 = (~(Wrxiu6 & Dsxiu6));
assign Dsxiu6 = (~(Qudpw6 & IRQ[12]));
assign Wrxiu6 = (Ksxiu6 & X6giu6);
assign X6giu6 = (~(Kwfiu6 & HWDATA[12]));
assign Ksxiu6 = (~(Odgpw6[12] & Rsxiu6));
assign Rsxiu6 = (~(K66iu6 & HWDATA[12]));
assign E7giu6 = (Sb5iu6 | Ysxiu6);
assign K2phu6 = (A5giu6 & Ftxiu6);
assign Ftxiu6 = (~(Mtxiu6 & Ttxiu6));
assign Ttxiu6 = (~(Vtdpw6 & IRQ[13]));
assign Mtxiu6 = (Auxiu6 & T4giu6);
assign T4giu6 = (~(Kwfiu6 & HWDATA[13]));
assign Auxiu6 = (~(Odgpw6[13] & Huxiu6));
assign Huxiu6 = (~(K66iu6 & HWDATA[13]));
assign A5giu6 = (Sb5iu6 | Ouxiu6);
assign D2phu6 = (W2giu6 & Vuxiu6);
assign Vuxiu6 = (~(Cvxiu6 & Jvxiu6));
assign Jvxiu6 = (~(Otdpw6 & IRQ[14]));
assign Cvxiu6 = (Qvxiu6 & P2giu6);
assign P2giu6 = (~(Kwfiu6 & HWDATA[14]));
assign Qvxiu6 = (~(Odgpw6[14] & Xvxiu6));
assign Xvxiu6 = (~(K66iu6 & HWDATA[14]));
assign W2giu6 = (~(Clfiu6 & R3giu6));
assign W1phu6 = (S0giu6 & Ewxiu6);
assign Ewxiu6 = (~(Lwxiu6 & Swxiu6));
assign Swxiu6 = (~(Lvdpw6 & IRQ[15]));
assign Lwxiu6 = (Zwxiu6 & L0giu6);
assign L0giu6 = (~(Fsdiu6 & Kwfiu6));
assign Zwxiu6 = (~(Odgpw6[15] & Gxxiu6));
assign Gxxiu6 = (~(Fsdiu6 & K66iu6));
assign Fsdiu6 = (Npdhu6 & HWDATA[15]);
assign S0giu6 = (Sb5iu6 | Nxxiu6);
assign P1phu6 = (Mvhiu6 & Uxxiu6);
assign Uxxiu6 = (~(Byxiu6 & Iyxiu6));
assign Iyxiu6 = (~(Atdpw6 & IRQ[16]));
assign Byxiu6 = (Pyxiu6 & Fvhiu6);
assign Fvhiu6 = (~(Kwfiu6 & HWDATA[16]));
assign Pyxiu6 = (~(Odgpw6[16] & Wyxiu6));
assign Wyxiu6 = (~(K66iu6 & HWDATA[16]));
assign Mvhiu6 = (~(Clfiu6 & Hwhiu6));
assign I1phu6 = (Npdiu6 & Dzxiu6);
assign Dzxiu6 = (~(Kzxiu6 & Rzxiu6));
assign Rzxiu6 = (~(Htdpw6 & IRQ[17]));
assign Kzxiu6 = (Yzxiu6 & Gpdiu6);
assign Gpdiu6 = (~(Kwfiu6 & HWDATA[17]));
assign Yzxiu6 = (~(Odgpw6[17] & F0yiu6));
assign F0yiu6 = (~(K66iu6 & HWDATA[17]));
assign Npdiu6 = (Sb5iu6 | M0yiu6);
assign B1phu6 = (Omdiu6 & T0yiu6);
assign T0yiu6 = (~(A1yiu6 & H1yiu6));
assign H1yiu6 = (~(Tsdpw6 & IRQ[18]));
assign A1yiu6 = (O1yiu6 & Hmdiu6);
assign Hmdiu6 = (~(Kwfiu6 & HWDATA[18]));
assign O1yiu6 = (~(Odgpw6[18] & V1yiu6));
assign V1yiu6 = (~(K66iu6 & HWDATA[18]));
assign Omdiu6 = (Sb5iu6 | C2yiu6);
assign U0phu6 = (Pjdiu6 & J2yiu6);
assign J2yiu6 = (~(Q2yiu6 & X2yiu6));
assign X2yiu6 = (~(Msdpw6 & IRQ[19]));
assign Q2yiu6 = (E3yiu6 & Ijdiu6);
assign Ijdiu6 = (~(Kwfiu6 & HWDATA[19]));
assign E3yiu6 = (~(Odgpw6[19] & L3yiu6));
assign L3yiu6 = (~(K66iu6 & HWDATA[19]));
assign Pjdiu6 = (Sb5iu6 | S3yiu6);
assign N0phu6 = (Qgdiu6 & Z3yiu6);
assign Z3yiu6 = (~(G4yiu6 & N4yiu6));
assign N4yiu6 = (~(Yrdpw6 & IRQ[20]));
assign G4yiu6 = (U4yiu6 & Jgdiu6);
assign Jgdiu6 = (~(Kwfiu6 & HWDATA[20]));
assign U4yiu6 = (~(Odgpw6[20] & B5yiu6));
assign B5yiu6 = (~(K66iu6 & HWDATA[20]));
assign Qgdiu6 = (Sb5iu6 | I5yiu6);
assign I5yiu6 = (!Lhdiu6);
assign G0phu6 = (Rddiu6 & P5yiu6);
assign P5yiu6 = (~(W5yiu6 & D6yiu6));
assign D6yiu6 = (~(Rrdpw6 & IRQ[21]));
assign W5yiu6 = (K6yiu6 & Kddiu6);
assign Kddiu6 = (~(Kwfiu6 & HWDATA[21]));
assign K6yiu6 = (~(Odgpw6[21] & R6yiu6));
assign R6yiu6 = (~(K66iu6 & HWDATA[21]));
assign Rddiu6 = (Sb5iu6 | Y6yiu6);
assign Zzohu6 = (Sadiu6 & F7yiu6);
assign F7yiu6 = (~(M7yiu6 & T7yiu6));
assign T7yiu6 = (~(Xndpw6 & IRQ[22]));
assign M7yiu6 = (A8yiu6 & Ladiu6);
assign Ladiu6 = (~(Kwfiu6 & HWDATA[22]));
assign A8yiu6 = (~(Odgpw6[22] & H8yiu6));
assign H8yiu6 = (~(K66iu6 & HWDATA[22]));
assign Sadiu6 = (Sb5iu6 | O8yiu6);
assign Szohu6 = (T7diu6 & V8yiu6);
assign V8yiu6 = (~(C9yiu6 & J9yiu6));
assign J9yiu6 = (~(Drdpw6 & IRQ[23]));
assign C9yiu6 = (Q9yiu6 & M7diu6);
assign M7diu6 = (~(Kwfiu6 & HWDATA[23]));
assign Q9yiu6 = (~(Odgpw6[23] & X9yiu6));
assign X9yiu6 = (~(K66iu6 & HWDATA[23]));
assign T7diu6 = (Sb5iu6 | Eayiu6);
assign Lzohu6 = (Nufiu6 & Layiu6);
assign Layiu6 = (~(Sayiu6 & Zayiu6));
assign Zayiu6 = (~(Pqdpw6 & IRQ[26]));
assign Sayiu6 = (Gbyiu6 & Gufiu6);
assign Gufiu6 = (~(Kwfiu6 & HWDATA[26]));
assign Gbyiu6 = (~(Odgpw6[26] & Nbyiu6));
assign Nbyiu6 = (~(K66iu6 & HWDATA[26]));
assign Nufiu6 = (Sb5iu6 | Ubyiu6);
assign Ezohu6 = (Jsfiu6 & Bcyiu6);
assign Bcyiu6 = (~(Icyiu6 & Pcyiu6));
assign Pcyiu6 = (~(Iqdpw6 & IRQ[27]));
assign Icyiu6 = (Wcyiu6 & Csfiu6);
assign Csfiu6 = (~(Kwfiu6 & HWDATA[27]));
assign Wcyiu6 = (~(Odgpw6[27] & Ddyiu6));
assign Ddyiu6 = (~(K66iu6 & HWDATA[27]));
assign Jsfiu6 = (Sb5iu6 | Kdyiu6);
assign Xyohu6 = (Fqfiu6 & Rdyiu6);
assign Rdyiu6 = (~(Ydyiu6 & Feyiu6));
assign Feyiu6 = (~(Bqdpw6 & IRQ[28]));
assign Ydyiu6 = (Meyiu6 & Ypfiu6);
assign Ypfiu6 = (~(Kwfiu6 & HWDATA[28]));
assign Meyiu6 = (~(Odgpw6[28] & Teyiu6));
assign Teyiu6 = (~(K66iu6 & HWDATA[28]));
assign Fqfiu6 = (Sb5iu6 | Afyiu6);
assign Qyohu6 = (Fgbiu6 & Hfyiu6);
assign Hfyiu6 = (~(Ofyiu6 & Vfyiu6));
assign Vfyiu6 = (~(Updpw6 & IRQ[29]));
assign Ofyiu6 = (Cgyiu6 & Yfbiu6);
assign Yfbiu6 = (~(Kwfiu6 & HWDATA[29]));
assign Cgyiu6 = (~(Odgpw6[29] & Jgyiu6));
assign Jgyiu6 = (~(K66iu6 & HWDATA[29]));
assign Fgbiu6 = (Sb5iu6 | Qgyiu6);
assign Jyohu6 = (Qxhiu6 & Xgyiu6);
assign Xgyiu6 = (~(Ehyiu6 & Lhyiu6));
assign Lhyiu6 = (~(Zvdpw6 & IRQ[30]));
assign Ehyiu6 = (Shyiu6 & Jxhiu6);
assign Jxhiu6 = (~(Kwfiu6 & HWDATA[30]));
assign Shyiu6 = (~(Odgpw6[30] & Zhyiu6));
assign Zhyiu6 = (~(K66iu6 & HWDATA[30]));
assign Qxhiu6 = (Sb5iu6 | Giyiu6);
assign Cyohu6 = (Bebiu6 & Niyiu6);
assign Niyiu6 = (~(Uiyiu6 & Bjyiu6));
assign Bjyiu6 = (~(Npdpw6 & IRQ[31]));
assign Uiyiu6 = (Ijyiu6 & Udbiu6);
assign Udbiu6 = (~(Kwfiu6 & HWDATA[31]));
assign Kwfiu6 = (Pjyiu6 & Yzciu6);
assign Yzciu6 = (Wjyiu6 & Npdhu6);
assign Ijyiu6 = (~(Odgpw6[31] & Dkyiu6));
assign Dkyiu6 = (~(K66iu6 & HWDATA[31]));
assign K66iu6 = (Kkyiu6 & D5eiu6);
assign Kkyiu6 = (Pjyiu6 & Npdhu6);
assign Bebiu6 = (~(Clfiu6 & Webiu6));
assign Clfiu6 = (!Sb5iu6);
assign Sb5iu6 = (~(Rkyiu6 & Ykyiu6));
assign Ykyiu6 = (~(Xe8iu6 | Ae0iu6));
assign Rkyiu6 = (~(G7oiu6 | Nloiu6));
assign Vxohu6 = (O25iu6 ? X3fpw6[3] : Flyiu6);
assign Flyiu6 = (~(Mlyiu6 & Tlyiu6));
assign Tlyiu6 = (Amyiu6 & Hmyiu6);
assign Hmyiu6 = (~(Omyiu6 & S8fpw6[11]));
assign Amyiu6 = (Vmyiu6 & Cnyiu6);
assign Cnyiu6 = (~(Jnyiu6 & D7fpw6[10]));
assign Jnyiu6 = (D7fpw6[6] & Qnyiu6);
assign Qnyiu6 = (Xiiiu6 | Mtjiu6);
assign Vmyiu6 = (~(L45iu6 & Xnyiu6));
assign Xnyiu6 = (Eoyiu6 | Loyiu6);
assign Loyiu6 = (Soyiu6 & N55iu6);
assign Soyiu6 = (~(K9aiu6 | Zoyiu6));
assign Mlyiu6 = (Gpyiu6 & Npyiu6);
assign Npyiu6 = (~(A95iu6 & D7fpw6[3]));
assign Oxohu6 = (Upyiu6 & Bqyiu6);
assign Bqyiu6 = (~(Iqyiu6 & Pqyiu6));
assign Pqyiu6 = (Wqyiu6 & Dryiu6);
assign Dryiu6 = (Kryiu6 & Rryiu6);
assign Rryiu6 = (Yryiu6 & O4aiu6);
assign Kryiu6 = (Fsyiu6 & Uloiu6);
assign Fsyiu6 = (~(Msyiu6 & Y0jiu6));
assign Msyiu6 = (~(Sijiu6 | Cyfpw6[3]));
assign Wqyiu6 = (Tsyiu6 & Atyiu6);
assign Atyiu6 = (~(Htyiu6 & Otyiu6));
assign Otyiu6 = (~(Vtyiu6 & Cuyiu6));
assign Cuyiu6 = (~(Juyiu6 & Quyiu6));
assign Juyiu6 = (Xuyiu6 & A95iu6);
assign Vtyiu6 = (~(Evyiu6 | P0piu6));
assign Tsyiu6 = (Lvyiu6 & Svyiu6);
assign Svyiu6 = (~(Zvyiu6 & Ae0iu6));
assign Zvyiu6 = (D6kiu6 & Gwyiu6);
assign Lvyiu6 = (~(W8aiu6 & Nwyiu6));
assign Nwyiu6 = (~(Uwyiu6 & Bxyiu6));
assign Bxyiu6 = (~(Ixyiu6 & Cyfpw6[7]));
assign Ixyiu6 = (Cyfpw6[5] & Pxyiu6);
assign Uwyiu6 = (Lkaiu6 | Wxyiu6);
assign Iqyiu6 = (Dyyiu6 & Kyyiu6);
assign Kyyiu6 = (Ryyiu6 & Yyyiu6);
assign Yyyiu6 = (Fzyiu6 & Mzyiu6);
assign Mzyiu6 = (~(Tzyiu6 & Geaiu6));
assign Tzyiu6 = (~(A0ziu6 & H0ziu6));
assign H0ziu6 = (O0ziu6 & V0ziu6);
assign V0ziu6 = (~(C1ziu6 & J1ziu6));
assign C1ziu6 = (~(Q1ziu6 | X1ziu6));
assign O0ziu6 = (E2ziu6 & Gjjiu6);
assign Gjjiu6 = (~(L2ziu6 & S2ziu6));
assign L2ziu6 = (L45iu6 & K9aiu6);
assign A0ziu6 = (Z2ziu6 & G3ziu6);
assign G3ziu6 = (~(U4kiu6 & N3ziu6));
assign Z2ziu6 = (~(D1piu6 & Xzmiu6));
assign Fzyiu6 = (~(Imaiu6 & U3ziu6));
assign U3ziu6 = (~(B4ziu6 & I4ziu6));
assign I4ziu6 = (~(W0piu6 & P4ziu6));
assign P4ziu6 = (~(W4ziu6 & D5ziu6));
assign D5ziu6 = (~(K5ziu6 & R5ziu6));
assign R5ziu6 = (~(Ndiiu6 ^ Y5ziu6));
assign K5ziu6 = (~(F6ziu6 | D7fpw6[13]));
assign W4ziu6 = (~(M6ziu6 & X1ziu6));
assign M6ziu6 = (~(T6ziu6 & A7ziu6));
assign A7ziu6 = (H7ziu6 & O7ziu6);
assign H7ziu6 = (~(V7ziu6 & C8ziu6));
assign C8ziu6 = (~(I6jiu6 | D7fpw6[4]));
assign V7ziu6 = (J8ziu6 & D7fpw6[11]);
assign T6ziu6 = (D7fpw6[13] & Q8ziu6);
assign Q8ziu6 = (~(X8ziu6 & Tniiu6));
assign B4ziu6 = (~(E9ziu6 & Q5aiu6));
assign E9ziu6 = (~(L9ziu6 & S9ziu6));
assign S9ziu6 = (~(Jiiiu6 & Z9ziu6));
assign Z9ziu6 = (~(Gaziu6 & Naziu6));
assign Naziu6 = (Oviiu6 | Gkiiu6);
assign L9ziu6 = (~(Dmiiu6 & Uaziu6));
assign Uaziu6 = (~(Bbziu6 & Ibziu6));
assign Ibziu6 = (~(D7fpw6[10] | D7fpw6[12]));
assign Bbziu6 = (Pbziu6 & Wbziu6);
assign Wbziu6 = (~(Dcziu6 ^ D7fpw6[9]));
assign Pbziu6 = (Ndiiu6 ? D7fpw6[7] : Kcziu6);
assign Ryyiu6 = (Rcziu6 & Ycziu6);
assign Ycziu6 = (E45iu6 | Wthiu6);
assign Dyyiu6 = (Fdziu6 & Mdziu6);
assign Mdziu6 = (D7fpw6[14] ? Aeziu6 : Tdziu6);
assign Aeziu6 = (~(Heziu6 & Nriiu6));
assign Heziu6 = (Aujiu6 & K9aiu6);
assign Fdziu6 = (Oeziu6 & Veziu6);
assign Upyiu6 = (H6ghu6 | HREADY);
assign Hxohu6 = (~(Cfziu6 & Jfziu6));
assign Jfziu6 = (Qfziu6 & Xfziu6);
assign Xfziu6 = (~(Egziu6 & Eafpw6[29]));
assign Qfziu6 = (Lgziu6 & Sgziu6);
assign Lgziu6 = (~(Zgziu6 & Fj8iu6));
assign Fj8iu6 = (~(Ghziu6 & Nhziu6));
assign Nhziu6 = (Uhziu6 & Biziu6);
assign Biziu6 = (Iiziu6 | Piziu6);
assign Uhziu6 = (Wiziu6 & Djziu6);
assign Wiziu6 = (Kjziu6 | Rjziu6);
assign Ghziu6 = (Yjziu6 & Fkziu6);
assign Fkziu6 = (Mkziu6 | Tkziu6);
assign Yjziu6 = (Alziu6 | Hlziu6);
assign Cfziu6 = (Olziu6 & Vlziu6);
assign Vlziu6 = (~(Zsfpw6[28] & Cmziu6));
assign Olziu6 = (~(vis_pc_o[28] & Jmziu6));
assign Axohu6 = (!Qmziu6);
assign Qmziu6 = (HREADY ? Xmziu6 : Tfjiu6);
assign Xmziu6 = (Enziu6 & Lnziu6);
assign Lnziu6 = (Snziu6 & Znziu6);
assign Znziu6 = (Goziu6 & Noziu6);
assign Noziu6 = (~(Bi0iu6 | Uoziu6));
assign Goziu6 = (Bpziu6 & Oaiiu6);
assign Bpziu6 = (~(Ipziu6 & Qe8iu6));
assign Snziu6 = (Ppziu6 & Wpziu6);
assign Wpziu6 = (~(Neoiu6 & Dqziu6));
assign Dqziu6 = (~(Kqziu6 & Rqziu6));
assign Rqziu6 = (~(Yqziu6 & D1piu6));
assign Yqziu6 = (Frziu6 & Cyfpw6[5]);
assign Kqziu6 = (Ntgiu6 & E4jiu6);
assign Ppziu6 = (Mrziu6 & Trziu6);
assign Trziu6 = (~(Asziu6 & Uriiu6));
assign Asziu6 = (~(Hsziu6 & Osziu6));
assign Osziu6 = (~(Vsziu6 & Ia8iu6));
assign Vsziu6 = (~(E4jiu6 | Cyfpw6[3]));
assign Hsziu6 = (Ctziu6 | Tfjiu6);
assign Mrziu6 = (Ctziu6 | As0iu6);
assign Enziu6 = (Jtziu6 & Qtziu6);
assign Qtziu6 = (Xtziu6 & Euziu6);
assign Euziu6 = (Luziu6 & Suziu6);
assign Suziu6 = (~(Cyfpw6[7] & Zuziu6));
assign Zuziu6 = (~(Gvziu6 & Nvziu6));
assign Nvziu6 = (Q5aiu6 | Uvziu6);
assign Gvziu6 = (Bwziu6 & Iwziu6);
assign Iwziu6 = (~(Pwziu6 & Wwziu6));
assign Pwziu6 = (~(Dxziu6 | Cyfpw6[0]));
assign Bwziu6 = (Jojiu6 | Ii0iu6);
assign Luziu6 = (~(Kxziu6 & Rxziu6));
assign Rxziu6 = (~(Yxziu6 & Fyziu6));
assign Fyziu6 = (Myziu6 & Tyziu6);
assign Tyziu6 = (~(Azziu6 & Hzziu6));
assign Azziu6 = (~(Tfjiu6 | D7fpw6[15]));
assign Myziu6 = (~(P0piu6 | Ozziu6));
assign Yxziu6 = (X3jiu6 & Vzziu6);
assign Vzziu6 = (~(U0aiu6 & D7fpw6[3]));
assign X3jiu6 = (Jjhiu6 | Uriiu6);
assign Xtziu6 = (Fniiu6 & C00ju6);
assign C00ju6 = (~(J00ju6 & Zraiu6));
assign J00ju6 = (~(Q00ju6 & X00ju6));
assign X00ju6 = (E10ju6 & L10ju6);
assign L10ju6 = (S10ju6 & Z10ju6);
assign Z10ju6 = (~(G20ju6 & N20ju6));
assign G20ju6 = (~(Nsaiu6 | Xe8iu6));
assign S10ju6 = (U20ju6 & W8oiu6);
assign U20ju6 = (~(B30ju6 & Mmjiu6));
assign B30ju6 = (I30ju6 & Gwyiu6);
assign E10ju6 = (P30ju6 & W30ju6);
assign W30ju6 = (~(Hzziu6 & D40ju6));
assign D40ju6 = (~(K40ju6 & R40ju6));
assign R40ju6 = (~(Y40ju6 & Ii0iu6));
assign K40ju6 = (F50ju6 & Xe8iu6);
assign F50ju6 = (~(M50ju6 & V9ghu6));
assign M50ju6 = (~(P0biu6 | Cyfpw6[6]));
assign P30ju6 = (T50ju6 & A60ju6);
assign A60ju6 = (~(Omyiu6 & H60ju6));
assign H60ju6 = (~(O60ju6 & V60ju6));
assign V60ju6 = (~(Wp0iu6 & Qyniu6));
assign T50ju6 = (~(Yljiu6 & C70ju6));
assign C70ju6 = (~(Cyfpw6[7] & J70ju6));
assign J70ju6 = (As0iu6 | Dxziu6);
assign Q00ju6 = (Q70ju6 & X70ju6);
assign X70ju6 = (E80ju6 & L80ju6);
assign L80ju6 = (S80ju6 | Ftjiu6);
assign E80ju6 = (Z80ju6 & G90ju6);
assign G90ju6 = (~(N90ju6 & Uriiu6));
assign N90ju6 = (~(U90ju6 & Ba0ju6));
assign Ba0ju6 = (Ia0ju6 & Pa0ju6);
assign Pa0ju6 = (~(Wa0ju6 & Db0ju6));
assign Wa0ju6 = (Nbkiu6 & Oviiu6);
assign Ia0ju6 = (Kb0ju6 & Rb0ju6);
assign U90ju6 = (Yb0ju6 & Fc0ju6);
assign Fc0ju6 = (~(P0piu6 & Mc0ju6));
assign Mc0ju6 = (~(Tc0ju6 & Ad0ju6));
assign Ad0ju6 = (Hd0ju6 & Od0ju6);
assign Hd0ju6 = (~(D7fpw6[8] & Vd0ju6));
assign Vd0ju6 = (U5jiu6 | Dcziu6);
assign Tc0ju6 = (Ce0ju6 & Je0ju6);
assign Ce0ju6 = (I6jiu6 ? Kcziu6 : Qe0ju6);
assign Yb0ju6 = (Xe0ju6 | H95iu6);
assign Z80ju6 = (~(J9kiu6 & Ef0ju6));
assign Ef0ju6 = (~(Lf0ju6 & Sf0ju6));
assign Sf0ju6 = (Zf0ju6 & Gg0ju6);
assign Gg0ju6 = (~(Ng0ju6 & Oviiu6));
assign Ng0ju6 = (~(I6jiu6 & Je0ju6));
assign Je0ju6 = (O95iu6 | D7fpw6[9]);
assign Zf0ju6 = (~(D7fpw6[13] & Ug0ju6));
assign Ug0ju6 = (~(Bh0ju6 & Ih0ju6));
assign Ih0ju6 = (Ph0ju6 | D7fpw6[4]);
assign Bh0ju6 = (Ndiiu6 | Wh0ju6);
assign Lf0ju6 = (Di0ju6 & Ki0ju6);
assign Ki0ju6 = (~(D7fpw6[12] & Ri0ju6));
assign Ri0ju6 = (~(Yi0ju6 & Fj0ju6));
assign Fj0ju6 = (Mj0ju6 & Tj0ju6);
assign Tj0ju6 = (~(Ak0ju6 & Zwciu6));
assign Mj0ju6 = (Hk0ju6 | Oviiu6);
assign Yi0ju6 = (Ok0ju6 & Vk0ju6);
assign Vk0ju6 = (Kcziu6 | D7fpw6[10]);
assign Ok0ju6 = (Ndiiu6 | Qxoiu6);
assign Di0ju6 = (Cl0ju6 | D7fpw6[7]);
assign Cl0ju6 = (!Zroiu6);
assign Q70ju6 = (~(Jl0ju6 | Ql0ju6));
assign Ql0ju6 = (~(Xl0ju6 | D7fpw6[8]));
assign Jl0ju6 = (C0ehu6 ? Lraiu6 : Em0ju6);
assign Em0ju6 = (Geoiu6 & H4ghu6);
assign Fniiu6 = (Hujiu6 | D7fpw6[12]);
assign Jtziu6 = (Lm0ju6 & F85iu6);
assign Lm0ju6 = (Sm0ju6 & Zm0ju6);
assign Zm0ju6 = (Wthiu6 | Nloiu6);
assign Sm0ju6 = (Taaiu6 | Faaiu6);
assign Twohu6 = (Gn0ju6 & Nn0ju6);
assign Nn0ju6 = (~(Un0ju6 & Bo0ju6));
assign Bo0ju6 = (Io0ju6 & Po0ju6);
assign Po0ju6 = (Wo0ju6 & Dp0ju6);
assign Dp0ju6 = (Kp0ju6 & Rp0ju6);
assign Rp0ju6 = (~(J9kiu6 & Yp0ju6));
assign Yp0ju6 = (~(Fq0ju6 & Mq0ju6));
assign Mq0ju6 = (Tq0ju6 & Ar0ju6);
assign Tq0ju6 = (~(D7fpw6[14] | D7fpw6[7]));
assign Fq0ju6 = (Hr0ju6 & D7fpw6[13]);
assign Hr0ju6 = (D7fpw6[5] & Or0ju6);
assign Or0ju6 = (~(Vr0ju6 & Cs0ju6));
assign Cs0ju6 = (~(Js0ju6 & Qs0ju6));
assign Qs0ju6 = (~(D7fpw6[4] | D7fpw6[6]));
assign Js0ju6 = (Wh0ju6 & F6ziu6);
assign Vr0ju6 = (~(Ak0ju6 & Oviiu6));
assign Kp0ju6 = (Xs0ju6 & Et0ju6);
assign Wo0ju6 = (Lt0ju6 & St0ju6);
assign St0ju6 = (~(Zt0ju6 & S6aiu6));
assign Zt0ju6 = (~(Ii0iu6 | Cyfpw6[4]));
assign Lt0ju6 = (~(Gu0ju6 & Xe8iu6));
assign Gu0ju6 = (W8aiu6 | M2piu6);
assign Io0ju6 = (Nu0ju6 & Uu0ju6);
assign Uu0ju6 = (Bv0ju6 & Iv0ju6);
assign Iv0ju6 = (~(Pv0ju6 & Mr0iu6));
assign Pv0ju6 = (Hzziu6 | N3ziu6);
assign Bv0ju6 = (~(Bziiu6 & D7fpw6[11]));
assign Nu0ju6 = (Wv0ju6 & Dw0ju6);
assign Dw0ju6 = (Kw0ju6 | Wxyiu6);
assign Wv0ju6 = (~(D7fpw6[14] & Rw0ju6));
assign Rw0ju6 = (~(Yw0ju6 & Fx0ju6));
assign Fx0ju6 = (Mx0ju6 & Tx0ju6);
assign Tx0ju6 = (~(Mtjiu6 & Ay0ju6));
assign Ay0ju6 = (~(Hy0ju6 & Oy0ju6));
assign Oy0ju6 = (Vy0ju6 & Oviiu6);
assign Vy0ju6 = (~(Cz0ju6 & Jz0ju6));
assign Cz0ju6 = (~(Hk0ju6 | D7fpw6[7]));
assign Hy0ju6 = (Qz0ju6 & Xz0ju6);
assign Xz0ju6 = (~(E01ju6 & D7fpw6[8]));
assign E01ju6 = (Tniiu6 ? L01ju6 : Dcziu6);
assign Mx0ju6 = (S01ju6 | Jjhiu6);
assign Yw0ju6 = (Z01ju6 & G11ju6);
assign G11ju6 = (Hk0ju6 | H95iu6);
assign Un0ju6 = (N11ju6 & U11ju6);
assign U11ju6 = (B21ju6 & I21ju6);
assign I21ju6 = (P21ju6 & W21ju6);
assign W21ju6 = (~(N3ziu6 & Taaiu6));
assign P21ju6 = (~(Y0jiu6 & D31ju6));
assign B21ju6 = (K31ju6 & R31ju6);
assign R31ju6 = (Nloiu6 | Lkaiu6);
assign K31ju6 = (Jjhiu6 | Y31ju6);
assign N11ju6 = (F41ju6 & M41ju6);
assign M41ju6 = (T41ju6 & A51ju6);
assign A51ju6 = (Wiliu6 | Ftjiu6);
assign F41ju6 = (~(H51ju6 | O51ju6));
assign O51ju6 = (Cyfpw6[6] ? V51ju6 : Yljiu6);
assign V51ju6 = (~(Ccoiu6 | R75iu6));
assign H51ju6 = (Cyfpw6[7] ? C61ju6 : M2piu6);
assign C61ju6 = (~(J61ju6 & Q61ju6));
assign Q61ju6 = (X61ju6 & E71ju6);
assign E71ju6 = (~(I30ju6 & Pxyiu6));
assign X61ju6 = (~(Moaiu6 & N2ghu6));
assign J61ju6 = (L71ju6 & S71ju6);
assign S71ju6 = (X5oiu6 | C0ehu6);
assign L71ju6 = (~(D1piu6 & Pugiu6));
assign Gn0ju6 = (Cyfpw6[7] | HREADY);
assign Mwohu6 = (G81ju6 ? H2fpw6[1] : Z71ju6);
assign Z71ju6 = (~(N81ju6 & U81ju6));
assign U81ju6 = (B91ju6 & I91ju6);
assign I91ju6 = (~(P91ju6 & D7fpw6[4]));
assign B91ju6 = (W91ju6 & Da1ju6);
assign Da1ju6 = (~(Ka1ju6 & Ra1ju6));
assign Ra1ju6 = (~(Jcaiu6 | D7fpw6[11]));
assign Ka1ju6 = (D7fpw6[13] & Ya1ju6);
assign W91ju6 = (~(Fb1ju6 & D7fpw6[9]));
assign N81ju6 = (Mb1ju6 & Tb1ju6);
assign Tb1ju6 = (~(D7fpw6[1] & Ac1ju6));
assign Fwohu6 = (Rgnhu6 & Hc1ju6);
assign Hc1ju6 = (~(Aw3iu6 & Oc1ju6));
assign Oc1ju6 = (~(Tonhu6 & Di1iu6));
assign Di1iu6 = (Tezhu6 & O8zhu6);
assign Tezhu6 = (Vc1ju6 & Cq3iu6);
assign Cq3iu6 = (Cd1ju6 & Fj1iu6);
assign Fj1iu6 = (Jd1ju6 & Qd1ju6);
assign Qd1ju6 = (Omzhu6 & Xj3iu6);
assign Xj3iu6 = (~(Xd1ju6 & Ow3iu6));
assign Ow3iu6 = (~(Ee1ju6 & Yn3iu6));
assign Yn3iu6 = (~(Ulnhu6 | Mdhpw6[2]));
assign Ee1ju6 = (Le1ju6 & Qnzhu6);
assign Qnzhu6 = (O8zhu6 | Mdhpw6[0]);
assign O8zhu6 = (!Mdhpw6[1]);
assign Le1ju6 = (~(Pinhu6 & Mdhpw6[1]));
assign Xd1ju6 = (~(Se1ju6 & Ze1ju6));
assign Ze1ju6 = (~(Fanhu6 | Jdnhu6));
assign Se1ju6 = (~(Ph1iu6 | Q8nhu6));
assign Ph1iu6 = (Gf1ju6 & X0ohu6);
assign Gf1ju6 = (Mo3iu6 & Aw3iu6);
assign Mo3iu6 = (Nf1ju6 & Uf1ju6);
assign Uf1ju6 = (~(Z63iu6 | Vmdpw6));
assign Z63iu6 = (G2ohu6 ^ Rrnhu6);
assign Nf1ju6 = (Rgnhu6 & Fmyhu6);
assign Fmyhu6 = (!N5yhu6);
assign N5yhu6 = (~(Bg1ju6 & Mdhpw6[3]));
assign Bg1ju6 = (U5yhu6 & Agyhu6);
assign Agyhu6 = (Ig1ju6 & Ighpw6[3]);
assign Ig1ju6 = (~(Vmzhu6 | Deyhu6));
assign Deyhu6 = (Zwyhu6 | Ighpw6[0]);
assign Zwyhu6 = (!Ighpw6[1]);
assign Omzhu6 = (~(Ighpw6[0] | Ighpw6[1]));
assign Jd1ju6 = (Iyyhu6 & U5yhu6);
assign Iyyhu6 = (Ez2iu6 & Wdyhu6);
assign Cd1ju6 = (~(Ulnhu6 | Mdhpw6[0]));
assign Vc1ju6 = (~(Vp3iu6 | Mdhpw6[2]));
assign Vp3iu6 = (~(Rzyhu6 ^ Mdhpw6[3]));
assign Rzyhu6 = (!Hknhu6);
assign Aw3iu6 = (!Yenhu6);
assign Yvohu6 = (Y14iu6 ? Mdhpw6[3] : Mdhpw6[2]);
assign Rvohu6 = (Y14iu6 ? Mdhpw6[2] : Mdhpw6[1]);
assign Y14iu6 = (!U03iu6);
assign Kvohu6 = (U03iu6 ? Mdhpw6[0] : Mdhpw6[1]);
assign Dvohu6 = (U03iu6 ? Ulnhu6 : Mdhpw6[0]);
assign U03iu6 = (Pg1ju6 & Wg1ju6);
assign Wg1ju6 = (~(Dh1ju6 & Ijzhu6));
assign Ijzhu6 = (~(Ighpw6[3] | Ighpw6[4]));
assign Dh1ju6 = (U5yhu6 & Vmzhu6);
assign Vmzhu6 = (!Ez2iu6);
assign Ez2iu6 = (Vuyhu6 & Eiyhu6);
assign Eiyhu6 = (!Ighpw6[4]);
assign Vuyhu6 = (!Ighpw6[2]);
assign Pg1ju6 = (~(Kh1ju6 & Rh1ju6));
assign Rh1ju6 = (Yh1ju6 & Pdyhu6);
assign Pdyhu6 = (!Pkyhu6);
assign Pkyhu6 = (Ighpw6[2] & Cvyhu6);
assign Yh1ju6 = (Cvyhu6 | Ighpw6[2]);
assign Cvyhu6 = (Ighpw6[0] & Ighpw6[1]);
assign Kh1ju6 = (Epyhu6 & U5yhu6);
assign U5yhu6 = (Vx2iu6 & Ujyhu6);
assign Vx2iu6 = (!Fnnhu6);
assign Epyhu6 = (Ighpw6[4] & Wdyhu6);
assign Wdyhu6 = (!Ighpw6[3]);
assign Wuohu6 = (O25iu6 ? X3fpw6[2] : Fi1ju6);
assign Fi1ju6 = (~(Mi1ju6 & Ti1ju6));
assign Ti1ju6 = (Aj1ju6 & Hj1ju6);
assign Hj1ju6 = (~(Omyiu6 & S8fpw6[10]));
assign Aj1ju6 = (Oj1ju6 & Vj1ju6);
assign Vj1ju6 = (~(D7fpw6[5] & K75iu6));
assign Oj1ju6 = (~(L45iu6 & N55iu6));
assign Mi1ju6 = (Ck1ju6 & Gpyiu6);
assign Ck1ju6 = (Jk1ju6 & Qk1ju6);
assign Qk1ju6 = (~(A95iu6 & D7fpw6[2]));
assign Jk1ju6 = (Ndiiu6 | H95iu6);
assign Puohu6 = (!Xk1ju6);
assign Xk1ju6 = (HREADY ? Ll1ju6 : El1ju6);
assign Ll1ju6 = (Sl1ju6 & Zl1ju6);
assign Iuohu6 = (!Gm1ju6);
assign Gm1ju6 = (HREADY ? Um1ju6 : Nm1ju6);
assign Um1ju6 = (Bn1ju6 & In1ju6);
assign In1ju6 = (Pn1ju6 & Wn1ju6);
assign Wn1ju6 = (Do1ju6 & Ko1ju6);
assign Ko1ju6 = (~(Ro1ju6 & Yo1ju6));
assign Ro1ju6 = (Fp1ju6 & Mp1ju6);
assign Mp1ju6 = (~(Ph0ju6 & Tp1ju6));
assign Tp1ju6 = (~(D7fpw6[7] & Aq1ju6));
assign Do1ju6 = (Hq1ju6 & Oq1ju6);
assign Pn1ju6 = (Vq1ju6 & Cr1ju6);
assign Cr1ju6 = (~(Oiaiu6 & Jr1ju6));
assign Jr1ju6 = (~(Qr1ju6 & Xr1ju6));
assign Xr1ju6 = (~(Es1ju6 & Qe8iu6));
assign Qr1ju6 = (~(Toaiu6 & Ls1ju6));
assign Vq1ju6 = (Ss1ju6 & Zs1ju6);
assign Zs1ju6 = (~(Gt1ju6 & M2piu6));
assign Gt1ju6 = (~(Ccoiu6 | Cyfpw6[0]));
assign Ss1ju6 = (~(K2aiu6 & Nt1ju6));
assign Nt1ju6 = (~(Ut1ju6 & Bu1ju6));
assign Bu1ju6 = (~(Iu1ju6 & Pu1ju6));
assign Iu1ju6 = (Md0iu6 & Sijiu6);
assign Ut1ju6 = (~(Qe8iu6 & Mr0iu6));
assign Bn1ju6 = (Wu1ju6 & Dv1ju6);
assign Dv1ju6 = (Kv1ju6 & Rv1ju6);
assign Rv1ju6 = (~(Yv1ju6 & Wliiu6));
assign Kv1ju6 = (Fw1ju6 & Mw1ju6);
assign Mw1ju6 = (~(Tw1ju6 & Oviiu6));
assign Tw1ju6 = (~(Ax1ju6 & Hx1ju6));
assign Hx1ju6 = (~(Yv1ju6 & Nbkiu6));
assign Fw1ju6 = (~(Pugiu6 & Ox1ju6));
assign Ox1ju6 = (~(Vx1ju6 & Cy1ju6));
assign Cy1ju6 = (~(M2piu6 & Jy1ju6));
assign Jy1ju6 = (~(Xojiu6 & Qy1ju6));
assign Qy1ju6 = (Mmjiu6 | Ae0iu6);
assign Wu1ju6 = (Xy1ju6 & Ez1ju6);
assign Xy1ju6 = (Lz1ju6 & Sz1ju6);
assign Sz1ju6 = (~(U98iu6 & Vxniu6));
assign Lz1ju6 = (Ax1ju6 | L01ju6);
assign Buohu6 = (~(Zz1ju6 & G02ju6));
assign G02ju6 = (~(C0ehu6 & N02ju6));
assign N02ju6 = (Eh6iu6 | Yv1ju6);
assign Zz1ju6 = (~(HREADY & U02ju6));
assign U02ju6 = (~(B12ju6 & I12ju6));
assign I12ju6 = (P12ju6 & W12ju6);
assign W12ju6 = (D22ju6 & K22ju6);
assign K22ju6 = (~(U98iu6 & R22ju6));
assign R22ju6 = (~(Y22ju6 & F32ju6));
assign F32ju6 = (M32ju6 | Xmliu6);
assign Y22ju6 = (~(Pthiu6 & Cyfpw6[1]));
assign D22ju6 = (T32ju6 & A42ju6);
assign T32ju6 = (~(H42ju6 & Neoiu6));
assign H42ju6 = (Omyiu6 & O42ju6);
assign O42ju6 = (~(V42ju6 & C52ju6));
assign C52ju6 = (J52ju6 & Q52ju6);
assign Q52ju6 = (As0iu6 | Xe8iu6);
assign J52ju6 = (X52ju6 & E62ju6);
assign X52ju6 = (L62ju6 | Cyfpw6[6]);
assign V42ju6 = (Cyfpw6[0] & S62ju6);
assign P12ju6 = (Z62ju6 & G72ju6);
assign G72ju6 = (~(Dxziu6 & N72ju6));
assign N72ju6 = (~(U72ju6 & B82ju6));
assign B82ju6 = (~(Ls1ju6 & Xzmiu6));
assign U72ju6 = (~(I82ju6 & Nlaiu6));
assign Z62ju6 = (P82ju6 | W82ju6);
assign B12ju6 = (D92ju6 & K92ju6);
assign K92ju6 = (R92ju6 & Y92ju6);
assign Y92ju6 = (~(Qe8iu6 & Fa2ju6));
assign Fa2ju6 = (~(Ma2ju6 & Ta2ju6));
assign Ta2ju6 = (H4ghu6 ? Hb2ju6 : Ab2ju6);
assign Hb2ju6 = (~(Dxziu6 & Ob2ju6));
assign Ob2ju6 = (~(Cyfpw6[5] & Vb2ju6));
assign Vb2ju6 = (~(Cc2ju6 & Eoyiu6));
assign Cc2ju6 = (~(Nlaiu6 | Cyfpw6[3]));
assign Ab2ju6 = (Jc2ju6 & Qc2ju6);
assign Qc2ju6 = (~(Xc2ju6 & Ed2ju6));
assign Ed2ju6 = (~(Xojiu6 | Sbghu6));
assign Xc2ju6 = (~(Nlaiu6 | Lkaiu6));
assign Ma2ju6 = (Ld2ju6 & M32ju6);
assign Ld2ju6 = (~(Sd2ju6 & Hs0iu6));
assign Sd2ju6 = (~(Q5aiu6 & Zd2ju6));
assign Zd2ju6 = (~(Fsdhu6 & Cqaiu6));
assign R92ju6 = (~(Yo1ju6 & I6jiu6));
assign D92ju6 = (Ge2ju6 & Ne2ju6);
assign Ne2ju6 = (~(W8aiu6 & Whfiu6));
assign Ge2ju6 = (D7fpw6[8] ? Bf2ju6 : Ue2ju6);
assign Bf2ju6 = (If2ju6 & Pf2ju6);
assign Pf2ju6 = (~(Wf2ju6 & Y5ziu6));
assign If2ju6 = (~(Yo1ju6 & Tniiu6));
assign Ue2ju6 = (Dg2ju6 & Kg2ju6);
assign Kg2ju6 = (~(Yo1ju6 & Rg2ju6));
assign Dg2ju6 = (Yg2ju6 & Fh2ju6);
assign Fh2ju6 = (~(Mh2ju6 & Htyiu6));
assign Mh2ju6 = (Th2ju6 & Ai2ju6);
assign Ai2ju6 = (~(Xe0ju6 & Hi2ju6));
assign Hi2ju6 = (~(Zroiu6 & Cwiiu6));
assign Yg2ju6 = (Oi2ju6 | Y5ziu6);
assign Y5ziu6 = (Vi2ju6 & Cj2ju6);
assign Cj2ju6 = (Jj2ju6 ^ Qj2ju6);
assign Qj2ju6 = (Xj2ju6 & Ek2ju6);
assign Ek2ju6 = (~(G8niu6 | Fp1ju6));
assign G8niu6 = (P9niu6 & vis_apsr_o[0]);
assign Xj2ju6 = (Lk2ju6 & Sk2ju6);
assign Sk2ju6 = (D7fpw6[11] | Qxoiu6);
assign Lk2ju6 = (Zk2ju6 | Gl2ju6);
assign Gl2ju6 = (Nl2ju6 ? Idfpw6[31] : Eafpw6[31]);
assign Zk2ju6 = (Ul2ju6 | P9niu6);
assign P9niu6 = (Bm2ju6 & Im2ju6);
assign Bm2ju6 = (Pm2ju6 & Wm2ju6);
assign Wm2ju6 = (~(Dn2ju6 & Kn2ju6));
assign Kn2ju6 = (~(Y2oiu6 | Tfjiu6));
assign Dn2ju6 = (~(Rn2ju6 | Yn2ju6));
assign Pm2ju6 = (~(Fo2ju6 & Mo2ju6));
assign Fo2ju6 = (~(Jjhiu6 | As0iu6));
assign Ul2ju6 = (~(Idfpw6[31] | Eafpw6[31]));
assign Idfpw6[31] = (To2ju6 & Oe0iu6);
assign Oe0iu6 = (~(Ap2ju6 & Hp2ju6));
assign Hp2ju6 = (Op2ju6 & Vp2ju6);
assign Vp2ju6 = (Cq2ju6 & Owaiu6);
assign Cq2ju6 = (~(Jq2ju6 & K9aiu6));
assign Jq2ju6 = (~(Knaiu6 & Qq2ju6));
assign Qq2ju6 = (Xe8iu6 | Cyfpw6[4]);
assign Op2ju6 = (Xq2ju6 & Er2ju6);
assign Er2ju6 = (Nlaiu6 | Lkaiu6);
assign Xq2ju6 = (~(F3aiu6 & Ldoiu6));
assign Ap2ju6 = (Lr2ju6 & Sr2ju6);
assign Sr2ju6 = (H6ghu6 & Zr2ju6);
assign Zr2ju6 = (~(Pthiu6 & H4ghu6));
assign Lr2ju6 = (~(Gs2ju6 | Ns2ju6));
assign Ns2ju6 = (Cyfpw6[4] ? Bt2ju6 : Us2ju6);
assign Bt2ju6 = (~(Wfoiu6 | R75iu6));
assign Gs2ju6 = (Cyfpw6[6] ? Pt2ju6 : It2ju6);
assign Jj2ju6 = (~(Wt2ju6 & Du2ju6));
assign Du2ju6 = (Fhoiu6 ? Ku2ju6 : Vioiu6);
assign Ku2ju6 = (!vis_apsr_o[3]);
assign Vioiu6 = (E5ehu6 ? Ru2ju6 : Bbliu6);
assign Wt2ju6 = (~(Fp1ju6 | Zroiu6));
assign Vi2ju6 = (Yu2ju6 & Fv2ju6);
assign Fv2ju6 = (Mv2ju6 | Tv2ju6);
assign Tv2ju6 = (Ng8iu6 ? vis_apsr_o[1] : Ri8iu6);
assign Ng8iu6 = (Aw2ju6 & Im2ju6);
assign Im2ju6 = (Hw2ju6 & Ow2ju6);
assign Ow2ju6 = (~(Vw2ju6 & Cx2ju6));
assign Cx2ju6 = (Jx2ju6 & Qx2ju6);
assign Qx2ju6 = (~(Xx2ju6 & Ey2ju6));
assign Xx2ju6 = (Mr0iu6 | Ly2ju6);
assign Jx2ju6 = (~(Sy2ju6 | Oiaiu6));
assign Vw2ju6 = (C0ehu6 & Zy2ju6);
assign Zy2ju6 = (Y2oiu6 | Qxaiu6);
assign Hw2ju6 = (~(Gz2ju6 | Nz2ju6));
assign Aw2ju6 = (Uz2ju6 & B03ju6);
assign B03ju6 = (~(C0ehu6 & I03ju6));
assign I03ju6 = (~(P03ju6 & O60ju6));
assign Uz2ju6 = (~(Cyfpw6[4] & W03ju6));
assign W03ju6 = (~(D13ju6 & K13ju6));
assign K13ju6 = (Mr0iu6 | Cyfpw6[7]);
assign D13ju6 = (R13ju6 & Y13ju6);
assign Y13ju6 = (~(F23ju6 & M23ju6));
assign M23ju6 = (Ii0iu6 | Pugiu6);
assign R13ju6 = (~(T23ju6 & Pfoiu6));
assign Ri8iu6 = (E5ehu6 ? A33ju6 : Caehu6);
assign A33ju6 = (~(H33ju6 & O33ju6));
assign O33ju6 = (~(V33ju6 & C43ju6));
assign C43ju6 = (J43ju6 & vis_apsr_o[1]);
assign V33ju6 = (~(Q43ju6 | X43ju6));
assign H33ju6 = (~(E53ju6 & L53ju6));
assign L53ju6 = (~(S53ju6 & Z53ju6));
assign S53ju6 = (~(X43ju6 | G63ju6));
assign E53ju6 = (~(N63ju6 & U63ju6));
assign U63ju6 = (~(B73ju6 & I73ju6));
assign I73ju6 = (~(P73ju6 & Cyfpw6[3]));
assign B73ju6 = (W73ju6 & Mr0iu6);
assign W73ju6 = (~(D83ju6 & K83ju6));
assign K83ju6 = (~(R83ju6 & Y83ju6));
assign R83ju6 = (~(F93ju6 | M93ju6));
assign D83ju6 = (~(T93ju6 & Aa3ju6));
assign Aa3ju6 = (~(Ha3ju6 & Oa3ju6));
assign T93ju6 = (F93ju6 ? Cb3ju6 : Va3ju6);
assign Cb3ju6 = (Jb3ju6 | Oa3ju6);
assign Va3ju6 = (Qb3ju6 & M93ju6);
assign N63ju6 = (P73ju6 ? Ru2ju6 : Xb3ju6);
assign P73ju6 = (Ec3ju6 & Q43ju6);
assign Ec3ju6 = (~(Lc3ju6 & Sc3ju6));
assign Lc3ju6 = (J43ju6 & Zc3ju6);
assign J43ju6 = (!G63ju6);
assign Ru2ju6 = (Gd3ju6 & Nd3ju6);
assign Nd3ju6 = (Ud3ju6 & Be3ju6);
assign Be3ju6 = (~(Ie3ju6 & Pe3ju6));
assign Ie3ju6 = (~(We3ju6 | Df3ju6));
assign Ud3ju6 = (Kf3ju6 | Ha3ju6);
assign Gd3ju6 = (~(Rf3ju6 | Yf3ju6));
assign Yf3ju6 = (~(Fg3ju6 | Mg3ju6));
assign Rf3ju6 = (Ah3ju6 ? Tg3ju6 : Jb3ju6);
assign Tg3ju6 = (Hh3ju6 & Oh3ju6);
assign Hh3ju6 = (Vh3ju6 & Fg3ju6);
assign Xb3ju6 = (~(H4ghu6 & Ci3ju6));
assign Ci3ju6 = (~(Ji3ju6 & Qi3ju6));
assign Qi3ju6 = (~(Xi3ju6 & Ej3ju6));
assign Xi3ju6 = (Lj3ju6 & M93ju6);
assign Ji3ju6 = (M93ju6 ? Zj3ju6 : Sj3ju6);
assign Zj3ju6 = (~(F93ju6 & Gk3ju6));
assign Sj3ju6 = (Ej3ju6 ? Uk3ju6 : Nk3ju6);
assign Mv2ju6 = (~(Bl3ju6 & I6jiu6));
assign Bl3ju6 = (Zroiu6 | Il3ju6);
assign Yu2ju6 = (~(Pl3ju6 & Wl3ju6));
assign Wl3ju6 = (Fp1ju6 | Il3ju6);
assign Pl3ju6 = (Xe0ju6 ^ Dm3ju6);
assign Dm3ju6 = (Fhoiu6 ? Km3ju6 : V7liu6);
assign Fhoiu6 = (Rm3ju6 & Mwniu6);
assign Mwniu6 = (Szniu6 | Yn2ju6);
assign Rm3ju6 = (~(C0ehu6 & Ym3ju6));
assign Ym3ju6 = (~(Fn3ju6 & Mn3ju6));
assign Mn3ju6 = (Tn3ju6 & Ao3ju6);
assign Ao3ju6 = (~(H4ghu6 & Ho3ju6));
assign Ho3ju6 = (~(Oo3ju6 & Vo3ju6));
assign Oo3ju6 = (~(Hs0iu6 | Cp3ju6));
assign Tn3ju6 = (Jp3ju6 & Qp3ju6);
assign Jp3ju6 = (~(Ly2ju6 & Cyfpw6[4]));
assign Fn3ju6 = (Xp3ju6 & Eq3ju6);
assign Eq3ju6 = (Ezniu6 | Cyfpw6[6]);
assign Xp3ju6 = (Lq3ju6 & P03ju6);
assign P03ju6 = (~(Sq3ju6 & Hs0iu6));
assign Lq3ju6 = (Ey2ju6 | As0iu6);
assign Km3ju6 = (!vis_apsr_o[2]);
assign V7liu6 = (E5ehu6 ? Gr3ju6 : Zq3ju6);
assign Gr3ju6 = (~(Nr3ju6 & Ur3ju6));
assign Ur3ju6 = (Bs3ju6 & Is3ju6);
assign Is3ju6 = (~(Ps3ju6 & Ws3ju6));
assign Ws3ju6 = (~(Dt3ju6 & Kt3ju6));
assign Kt3ju6 = (Rt3ju6 & Yt3ju6);
assign Rt3ju6 = (~(Lj3ju6 | Jb3ju6));
assign Dt3ju6 = (Fu3ju6 & Mu3ju6);
assign Fu3ju6 = (Hv3ju6 ? Av3ju6 : Tu3ju6);
assign Av3ju6 = (Ov3ju6 & Vv3ju6);
assign Vv3ju6 = (~(Cw3ju6 | Jw3ju6));
assign Tu3ju6 = (Qw3ju6 & Xw3ju6);
assign Xw3ju6 = (~(Ex3ju6 | Lx3ju6));
assign Qw3ju6 = (~(Sx3ju6 | Zx3ju6));
assign Ps3ju6 = (~(Gy3ju6 & Oh3ju6));
assign Gy3ju6 = (Ah3ju6 & Ny3ju6);
assign Bs3ju6 = (Uy3ju6 & Bz3ju6);
assign Uy3ju6 = (~(Iz3ju6 & Pz3ju6));
assign Pz3ju6 = (~(Wz3ju6 & D04ju6));
assign D04ju6 = (K04ju6 & R04ju6);
assign K04ju6 = (Ha3ju6 & Uk3ju6);
assign Wz3ju6 = (Y04ju6 & F14ju6);
assign Y04ju6 = (Hv3ju6 ? T14ju6 : M14ju6);
assign T14ju6 = (A24ju6 & H24ju6);
assign H24ju6 = (~(O24ju6 | V24ju6));
assign A24ju6 = (C34ju6 & J34ju6);
assign M14ju6 = (Q34ju6 & X34ju6);
assign X34ju6 = (~(E44ju6 | L44ju6));
assign Iz3ju6 = (~(S44ju6 & Kf3ju6));
assign S44ju6 = (Z44ju6 & Ny3ju6);
assign Nr3ju6 = (G54ju6 & N54ju6);
assign N54ju6 = (~(U54ju6 & B64ju6));
assign B64ju6 = (~(I64ju6 & P64ju6));
assign P64ju6 = (W64ju6 & D74ju6);
assign D74ju6 = (K74ju6 & R74ju6);
assign R74ju6 = (~(Hv3ju6 & Y74ju6));
assign Y74ju6 = (F84ju6 | M84ju6);
assign K74ju6 = (T84ju6 & A94ju6);
assign W64ju6 = (H94ju6 & O94ju6);
assign H94ju6 = (~(M84ju6 & V94ju6));
assign I64ju6 = (Ca4ju6 & Ja4ju6);
assign Ja4ju6 = (Mg3ju6 & Qa4ju6);
assign Qa4ju6 = (~(F84ju6 & O24ju6));
assign Ca4ju6 = (~(Xa4ju6 | Eb4ju6));
assign G54ju6 = (~(Lb4ju6 & Sb4ju6));
assign Sb4ju6 = (~(Zb4ju6 & Gc4ju6));
assign Gc4ju6 = (Nc4ju6 & Uc4ju6);
assign Nc4ju6 = (~(Gk3ju6 | Y83ju6));
assign Zb4ju6 = (Bd4ju6 & Id4ju6);
assign Bd4ju6 = (Hv3ju6 ? Wd4ju6 : Pd4ju6);
assign Wd4ju6 = (Q34ju6 & De4ju6);
assign De4ju6 = (~(Ke4ju6 | Re4ju6));
assign Q34ju6 = (~(Ye4ju6 | Ff4ju6));
assign Pd4ju6 = (Ov3ju6 & Mf4ju6);
assign Mf4ju6 = (~(Tf4ju6 | Ag4ju6));
assign Ov3ju6 = (~(Hg4ju6 | Og4ju6));
assign Lb4ju6 = (~(Vg4ju6 & Oh3ju6));
assign Vg4ju6 = (Ch4ju6 & Ny3ju6);
assign Zq3ju6 = (~(Jh4ju6 & Qh4ju6));
assign Qh4ju6 = (Xh4ju6 & Ei4ju6);
assign Ei4ju6 = (Li4ju6 & Si4ju6);
assign Si4ju6 = (Zi4ju6 & Gj4ju6);
assign Gj4ju6 = (Ibliu6 & Kkkiu6);
assign Kkkiu6 = (Nj4ju6 & Uj4ju6);
assign Uj4ju6 = (Bk4ju6 & Ik4ju6);
assign Ik4ju6 = (~(Pk4ju6 & vis_ipsr_o[4]));
assign Bk4ju6 = (~(Affpw6[4] | Wk4ju6));
assign Nj4ju6 = (Dl4ju6 & Kl4ju6);
assign Kl4ju6 = (Eg0iu6 ? Yl4ju6 : Rl4ju6);
assign Eg0iu6 = (Mm4ju6 ? Fm4ju6 : V3iiu6);
assign Fm4ju6 = (Tm4ju6 & An4ju6);
assign An4ju6 = (Hn4ju6 & On4ju6);
assign On4ju6 = (Vn4ju6 & Co4ju6);
assign Co4ju6 = (~(Jo4ju6 & vis_r14_o[4]));
assign Vn4ju6 = (Qo4ju6 & Xo4ju6);
assign Xo4ju6 = (~(Ep4ju6 & vis_psp_o[2]));
assign Qo4ju6 = (~(Lp4ju6 & vis_msp_o[2]));
assign Hn4ju6 = (Sp4ju6 & Zp4ju6);
assign Zp4ju6 = (~(Gq4ju6 & vis_r12_o[4]));
assign Sp4ju6 = (~(Nq4ju6 & vis_r11_o[4]));
assign Tm4ju6 = (Uq4ju6 & Br4ju6);
assign Br4ju6 = (Ir4ju6 & Pr4ju6);
assign Pr4ju6 = (~(Wr4ju6 & vis_r10_o[4]));
assign Ir4ju6 = (~(Ds4ju6 & vis_r9_o[4]));
assign Uq4ju6 = (D50iu6 & Ks4ju6);
assign Ks4ju6 = (~(Rs4ju6 & vis_r8_o[4]));
assign V3iiu6 = (!Fkfpw6[4]);
assign Yl4ju6 = (~(Ys4ju6 & Qbfpw6[4]));
assign Rl4ju6 = (~(Ft4ju6 | Mt4ju6));
assign Ft4ju6 = (Qbfpw6[4] ? Tt4ju6 : Ys4ju6);
assign Qbfpw6[4] = (~(Au4ju6 ^ Hu4ju6));
assign Au4ju6 = (~(Ou4ju6 & Vu4ju6));
assign Vu4ju6 = (Cv4ju6 & Jv4ju6);
assign Jv4ju6 = (B5kiu6 | Qv4ju6);
assign Cv4ju6 = (~(S8fpw6[4] & Xv4ju6));
assign Ou4ju6 = (Ew4ju6 & Lw4ju6);
assign Lw4ju6 = (~(Sw4ju6 & Zw4ju6));
assign Ew4ju6 = (V4aiu6 | Gx4ju6);
assign Dl4ju6 = (Nx4ju6 & Ux4ju6);
assign Ux4ju6 = (~(By4ju6 & Eafpw6[4]));
assign Nx4ju6 = (~(Iy4ju6 & Zw4ju6));
assign Ibliu6 = (Py4ju6 & Wy4ju6);
assign Wy4ju6 = (Dz4ju6 & Kz4ju6);
assign Kz4ju6 = (~(Affpw6[0] | Wk4ju6));
assign Dz4ju6 = (Rz4ju6 & Yz4ju6);
assign Yz4ju6 = (~(F05ju6 & M05ju6));
assign M05ju6 = (~(Qjoiu6 | S8fpw6[2]));
assign F05ju6 = (T05ju6 & vis_primask_o);
assign Rz4ju6 = (~(Pk4ju6 & vis_ipsr_o[0]));
assign Py4ju6 = (A15ju6 & H15ju6);
assign H15ju6 = (Go0iu6 ? V15ju6 : O15ju6);
assign V15ju6 = (~(C25ju6 | Mt4ju6));
assign C25ju6 = (Qbfpw6[0] ? Tt4ju6 : Ys4ju6);
assign O15ju6 = (~(Ys4ju6 & Qbfpw6[0]));
assign Qbfpw6[0] = (~(J25ju6 ^ Hu4ju6));
assign J25ju6 = (~(Q25ju6 & X25ju6));
assign X25ju6 = (~(S8fpw6[0] & E35ju6));
assign Q25ju6 = (~(Sw4ju6 & L35ju6));
assign A15ju6 = (S35ju6 & Z35ju6);
assign Z35ju6 = (~(By4ju6 & Eafpw6[0]));
assign S35ju6 = (~(Iy4ju6 & L35ju6));
assign Zi4ju6 = (K5liu6 & Bbliu6);
assign Bbliu6 = (G45ju6 & N45ju6);
assign N45ju6 = (U45ju6 & B55ju6);
assign B55ju6 = (~(vis_apsr_o[3] & I55ju6));
assign U45ju6 = (~(Affpw6[31] | Wk4ju6));
assign G45ju6 = (P55ju6 & W55ju6);
assign W55ju6 = (To2ju6 ? K65ju6 : D65ju6);
assign To2ju6 = (!R65ju6);
assign K65ju6 = (~(Y65ju6 | Mt4ju6));
assign Y65ju6 = (Nl2ju6 ? Ys4ju6 : Tt4ju6);
assign Nl2ju6 = (!D5epw6);
assign D65ju6 = (~(Ys4ju6 & D5epw6));
assign D5epw6 = (F75ju6 | M75ju6);
assign F75ju6 = (Aioiu6 ? A85ju6 : T75ju6);
assign P55ju6 = (H85ju6 & O85ju6);
assign O85ju6 = (~(By4ju6 & Eafpw6[31]));
assign H85ju6 = (~(Iy4ju6 & Aioiu6));
assign K5liu6 = (V85ju6 & C95ju6);
assign C95ju6 = (J95ju6 & Q95ju6);
assign Q95ju6 = (~(X95ju6 & Sg0iu6));
assign X95ju6 = (Ys4ju6 & Qbfpw6[30]);
assign J95ju6 = (~(Affpw6[30] | Ea5ju6));
assign Ea5ju6 = (Iy4ju6 & T6liu6);
assign V85ju6 = (La5ju6 & Sa5ju6);
assign Sa5ju6 = (~(Za5ju6 & Gb5ju6));
assign Gb5ju6 = (Nb5ju6 | Ub5ju6);
assign Nb5ju6 = (Mt4ju6 | Qbfpw6[30]);
assign Za5ju6 = (~(Bc5ju6 & Ic5ju6));
assign Bc5ju6 = (Sg0iu6 | Pc5ju6);
assign Pc5ju6 = (Wc5ju6 & Qbfpw6[30]);
assign Qbfpw6[30] = (Dd5ju6 | M75ju6);
assign Dd5ju6 = (T6liu6 ? A85ju6 : T75ju6);
assign La5ju6 = (Kd5ju6 & Rd5ju6);
assign Rd5ju6 = (~(vis_apsr_o[2] & I55ju6));
assign Kd5ju6 = (~(By4ju6 & Eafpw6[30]));
assign Li4ju6 = (Yd5ju6 & Fe5ju6);
assign Fe5ju6 = (Cgkiu6 & Evkiu6);
assign Evkiu6 = (Me5ju6 & Te5ju6);
assign Te5ju6 = (Af5ju6 & Hf5ju6);
assign Hf5ju6 = (~(By4ju6 & Eafpw6[23]));
assign Af5ju6 = (~(Affpw6[23] | Of5ju6));
assign Of5ju6 = (~(Vf5ju6 | Fk0iu6));
assign Vf5ju6 = (Qbfpw6[23] ? Wc5ju6 : Cg5ju6);
assign Me5ju6 = (Jg5ju6 & Qg5ju6);
assign Qg5ju6 = (~(Iy4ju6 & Xg5ju6));
assign Jg5ju6 = (~(Ub5ju6 & Eh5ju6));
assign Eh5ju6 = (~(Lh5ju6 & Ic5ju6));
assign Lh5ju6 = (~(Fk0iu6 & Qbfpw6[23]));
assign Qbfpw6[23] = (~(Sh5ju6 ^ Hu4ju6));
assign Sh5ju6 = (Zh5ju6 | Gi5ju6);
assign Gi5ju6 = (D7fpw6[13] ? Ui5ju6 : Ni5ju6);
assign Ni5ju6 = (~(Gx4ju6 | S8fpw6[11]));
assign Zh5ju6 = (~(Bj5ju6 & Ij5ju6));
assign Bj5ju6 = (~(Sw4ju6 & Xg5ju6));
assign Cgkiu6 = (Pj5ju6 & Wj5ju6);
assign Wj5ju6 = (Dk5ju6 & Kk5ju6);
assign Kk5ju6 = (~(Affpw6[2] | Rk5ju6));
assign Rk5ju6 = (Yk5ju6 & L8ehu6);
assign Yk5ju6 = (P8oiu6 & H6ghu6);
assign Dk5ju6 = (Fl5ju6 & Ml5ju6);
assign Ml5ju6 = (~(Pk4ju6 & vis_ipsr_o[2]));
assign Fl5ju6 = (~(By4ju6 & Eafpw6[2]));
assign Pj5ju6 = (Tl5ju6 & Am5ju6);
assign Am5ju6 = (Gh0iu6 ? Om5ju6 : Hm5ju6);
assign Gh0iu6 = (Cn5ju6 ? Fkfpw6[2] : Vm5ju6);
assign Vm5ju6 = (~(Jn5ju6 & Qn5ju6));
assign Qn5ju6 = (Xn5ju6 & Eo5ju6);
assign Eo5ju6 = (Lo5ju6 & So5ju6);
assign So5ju6 = (~(Jo4ju6 & vis_r14_o[2]));
assign Lo5ju6 = (Zo5ju6 & Gp5ju6);
assign Gp5ju6 = (~(Ep4ju6 & vis_psp_o[0]));
assign Zo5ju6 = (~(Lp4ju6 & vis_msp_o[0]));
assign Xn5ju6 = (Np5ju6 & Up5ju6);
assign Up5ju6 = (~(Gq4ju6 & vis_r12_o[2]));
assign Np5ju6 = (~(Nq4ju6 & vis_r11_o[2]));
assign Jn5ju6 = (Bq5ju6 & Iq5ju6);
assign Iq5ju6 = (Pq5ju6 & Wq5ju6);
assign Wq5ju6 = (~(Wr4ju6 & vis_r10_o[2]));
assign Pq5ju6 = (~(Ds4ju6 & vis_r9_o[2]));
assign Bq5ju6 = (F60iu6 & Dr5ju6);
assign Dr5ju6 = (~(Rs4ju6 & vis_r8_o[2]));
assign Om5ju6 = (~(Kr5ju6 | Mt4ju6));
assign Kr5ju6 = (Qbfpw6[2] ? Tt4ju6 : Ys4ju6);
assign Hm5ju6 = (~(Ys4ju6 & Qbfpw6[2]));
assign Qbfpw6[2] = (~(Rr5ju6 ^ Hu4ju6));
assign Rr5ju6 = (~(Yr5ju6 & Fs5ju6));
assign Fs5ju6 = (Ms5ju6 & Ts5ju6);
assign Ts5ju6 = (~(S8fpw6[2] & E35ju6));
assign Ms5ju6 = (Je8iu6 | Qv4ju6);
assign Yr5ju6 = (At5ju6 & Ht5ju6);
assign Ht5ju6 = (~(Sw4ju6 & Ot5ju6));
assign At5ju6 = (Ccaiu6 | Gx4ju6);
assign Tl5ju6 = (Vt5ju6 & Cu5ju6);
assign Cu5ju6 = (~(Iy4ju6 & Ot5ju6));
assign Vt5ju6 = (~(vis_control_o & Wk4ju6));
assign Yd5ju6 = (Lokiu6 & Dkkiu6);
assign Dkkiu6 = (Ju5ju6 & Qu5ju6);
assign Qu5ju6 = (Xu5ju6 & Ev5ju6);
assign Ev5ju6 = (~(By4ju6 & Eafpw6[3]));
assign Xu5ju6 = (~(Affpw6[3] | Lv5ju6));
assign Lv5ju6 = (Pk4ju6 & vis_ipsr_o[3]);
assign Ju5ju6 = (Sv5ju6 & Zv5ju6);
assign Zv5ju6 = (Lg0iu6 ? Nw5ju6 : Gw5ju6);
assign Lg0iu6 = (Mm4ju6 ? Uw5ju6 : Wjkiu6);
assign Uw5ju6 = (Bx5ju6 & Ix5ju6);
assign Ix5ju6 = (Px5ju6 & Wx5ju6);
assign Wx5ju6 = (Dy5ju6 & Ky5ju6);
assign Ky5ju6 = (~(Jo4ju6 & vis_r14_o[3]));
assign Dy5ju6 = (Ry5ju6 & Yy5ju6);
assign Yy5ju6 = (~(Ep4ju6 & vis_psp_o[1]));
assign Ry5ju6 = (~(Lp4ju6 & vis_msp_o[1]));
assign Px5ju6 = (Fz5ju6 & Mz5ju6);
assign Mz5ju6 = (~(Gq4ju6 & vis_r12_o[3]));
assign Fz5ju6 = (~(Nq4ju6 & vis_r11_o[3]));
assign Bx5ju6 = (Tz5ju6 & A06ju6);
assign A06ju6 = (H06ju6 & O06ju6);
assign O06ju6 = (~(Wr4ju6 & vis_r10_o[3]));
assign H06ju6 = (~(Ds4ju6 & vis_r9_o[3]));
assign Tz5ju6 = (K50iu6 & V06ju6);
assign V06ju6 = (~(Rs4ju6 & vis_r8_o[3]));
assign Wjkiu6 = (!Fkfpw6[3]);
assign Nw5ju6 = (~(Ys4ju6 & Qbfpw6[3]));
assign Gw5ju6 = (~(C16ju6 | Mt4ju6));
assign C16ju6 = (Qbfpw6[3] ? Tt4ju6 : Ys4ju6);
assign Qbfpw6[3] = (~(J16ju6 ^ Hu4ju6));
assign J16ju6 = (~(Q16ju6 & X16ju6));
assign X16ju6 = (E26ju6 & L26ju6);
assign L26ju6 = (Y8biu6 | Qv4ju6);
assign E26ju6 = (~(S8fpw6[3] & Xv4ju6));
assign Q16ju6 = (S26ju6 & Z26ju6);
assign Z26ju6 = (~(Sw4ju6 & G36ju6));
assign S26ju6 = (Prjiu6 | Gx4ju6);
assign Sv5ju6 = (N36ju6 & U36ju6);
assign U36ju6 = (~(Iy4ju6 & G36ju6));
assign N36ju6 = (~(Hlliu6 & Wk4ju6));
assign Lokiu6 = (B46ju6 & I46ju6);
assign I46ju6 = (P46ju6 & W46ju6);
assign W46ju6 = (~(Pk4ju6 & vis_ipsr_o[5]));
assign P46ju6 = (~(Affpw6[5] | Wk4ju6));
assign B46ju6 = (D56ju6 & K56ju6);
assign K56ju6 = (Xf0iu6 ? Y56ju6 : R56ju6);
assign Xf0iu6 = (Mm4ju6 ? F66ju6 : Eokiu6);
assign F66ju6 = (M66ju6 & T66ju6);
assign T66ju6 = (A76ju6 & H76ju6);
assign H76ju6 = (O76ju6 & V76ju6);
assign V76ju6 = (~(Jo4ju6 & vis_r14_o[5]));
assign O76ju6 = (C86ju6 & J86ju6);
assign J86ju6 = (~(Ep4ju6 & vis_psp_o[3]));
assign C86ju6 = (~(Lp4ju6 & vis_msp_o[3]));
assign A76ju6 = (Q86ju6 & X86ju6);
assign X86ju6 = (~(Gq4ju6 & vis_r12_o[5]));
assign Q86ju6 = (~(Nq4ju6 & vis_r11_o[5]));
assign M66ju6 = (E96ju6 & L96ju6);
assign L96ju6 = (S96ju6 & Z96ju6);
assign Z96ju6 = (~(Wr4ju6 & vis_r10_o[5]));
assign S96ju6 = (~(Ds4ju6 & vis_r9_o[5]));
assign E96ju6 = (W40iu6 & Ga6ju6);
assign Ga6ju6 = (~(Rs4ju6 & vis_r8_o[5]));
assign Eokiu6 = (!Fkfpw6[5]);
assign Y56ju6 = (~(Ys4ju6 & Qbfpw6[5]));
assign R56ju6 = (~(Na6ju6 | Mt4ju6));
assign Na6ju6 = (Qbfpw6[5] ? Tt4ju6 : Ys4ju6);
assign Qbfpw6[5] = (~(Ua6ju6 ^ Hu4ju6));
assign Ua6ju6 = (~(Bb6ju6 & Ib6ju6));
assign Ib6ju6 = (Pb6ju6 & Wb6ju6);
assign Wb6ju6 = (Cajiu6 | Qv4ju6);
assign Qv4ju6 = (~(Dc6ju6 | Kc6ju6));
assign Dc6ju6 = (H6ghu6 & Rc6ju6);
assign Rc6ju6 = (~(Yc6ju6 & Fd6ju6));
assign Fd6ju6 = (Md6ju6 & Fmjiu6);
assign Md6ju6 = (~(Td6ju6 & Cyfpw6[7]));
assign Td6ju6 = (Ae6ju6 & Jjhiu6);
assign Ae6ju6 = (~(He6ju6 & Oe6ju6));
assign Oe6ju6 = (X5oiu6 | Tfjiu6);
assign Yc6ju6 = (Ve6ju6 & Cf6ju6);
assign Cf6ju6 = (~(Cyfpw6[0] & F1jiu6));
assign F1jiu6 = (Xzmiu6 | Toaiu6);
assign Ve6ju6 = (~(Jf6ju6 & Oiaiu6));
assign Pb6ju6 = (~(S8fpw6[5] & Xv4ju6));
assign Bb6ju6 = (Qf6ju6 & Xf6ju6);
assign Xf6ju6 = (~(Sw4ju6 & Eg6ju6));
assign Qf6ju6 = (Gx4ju6 | A1kiu6);
assign D56ju6 = (Lg6ju6 & Sg6ju6);
assign Sg6ju6 = (~(By4ju6 & Eafpw6[5]));
assign Lg6ju6 = (~(Iy4ju6 & Eg6ju6));
assign Xh4ju6 = (Zg6ju6 & Gh6ju6);
assign Gh6ju6 = (Nh6ju6 & Uh6ju6);
assign Uh6ju6 = (~(Jukiu6 | Pqkiu6));
assign Pqkiu6 = (~(Bi6ju6 & Ii6ju6));
assign Ii6ju6 = (Pi6ju6 & Wi6ju6);
assign Wi6ju6 = (~(By4ju6 & Eafpw6[6]));
assign Pi6ju6 = (~(Affpw6[6] | Dj6ju6));
assign Dj6ju6 = (Iy4ju6 & Kj6ju6);
assign Bi6ju6 = (Rj6ju6 & Yj6ju6);
assign Yj6ju6 = (Fk6ju6 | Mk6ju6);
assign Fk6ju6 = (E2epw6 ? Wc5ju6 : Cg5ju6);
assign Rj6ju6 = (~(Ub5ju6 & Tk6ju6));
assign Tk6ju6 = (~(Al6ju6 & Ic5ju6));
assign Al6ju6 = (~(Mk6ju6 & E2epw6));
assign E2epw6 = (Hl6ju6 ^ Ol6ju6);
assign Hl6ju6 = (~(Vl6ju6 & Cm6ju6));
assign Cm6ju6 = (Jm6ju6 & Qm6ju6);
assign Qm6ju6 = (~(Kc6ju6 & S8fpw6[4]));
assign Jm6ju6 = (~(S8fpw6[6] & Xv4ju6));
assign Vl6ju6 = (Xm6ju6 & En6ju6);
assign En6ju6 = (~(Sw4ju6 & Kj6ju6));
assign Xm6ju6 = (Gx4ju6 | Dzjiu6);
assign Mk6ju6 = (!Qf0iu6);
assign Jukiu6 = (~(Ln6ju6 & Sn6ju6));
assign Sn6ju6 = (Zn6ju6 & Go6ju6);
assign Go6ju6 = (~(By4ju6 & Eafpw6[7]));
assign Zn6ju6 = (~(Affpw6[7] | No6ju6));
assign No6ju6 = (Iy4ju6 & Uo6ju6);
assign Ln6ju6 = (Bp6ju6 & Ip6ju6);
assign Ip6ju6 = (~(Ub5ju6 & Pp6ju6));
assign Pp6ju6 = (~(Wp6ju6 & Ic5ju6));
assign Wp6ju6 = (~(Jf0iu6 & S2epw6));
assign Bp6ju6 = (Dq6ju6 | Jf0iu6);
assign Jf0iu6 = (Mm4ju6 ? Kq6ju6 : Cukiu6);
assign Kq6ju6 = (Rq6ju6 & Yq6ju6);
assign Yq6ju6 = (Fr6ju6 & Mr6ju6);
assign Mr6ju6 = (Tr6ju6 & As6ju6);
assign As6ju6 = (~(Jo4ju6 & vis_r14_o[7]));
assign Tr6ju6 = (Hs6ju6 & Os6ju6);
assign Os6ju6 = (~(Ep4ju6 & vis_psp_o[5]));
assign Hs6ju6 = (~(Lp4ju6 & vis_msp_o[5]));
assign Fr6ju6 = (Vs6ju6 & Ct6ju6);
assign Ct6ju6 = (~(Gq4ju6 & vis_r12_o[7]));
assign Vs6ju6 = (~(Nq4ju6 & vis_r11_o[7]));
assign Rq6ju6 = (Jt6ju6 & Qt6ju6);
assign Qt6ju6 = (Xt6ju6 & Eu6ju6);
assign Eu6ju6 = (~(Wr4ju6 & vis_r10_o[7]));
assign Xt6ju6 = (~(Ds4ju6 & vis_r9_o[7]));
assign Jt6ju6 = (I40iu6 & Lu6ju6);
assign Lu6ju6 = (~(Rs4ju6 & vis_r8_o[7]));
assign Cukiu6 = (!Fkfpw6[7]);
assign Dq6ju6 = (S2epw6 ? Wc5ju6 : Cg5ju6);
assign S2epw6 = (~(Su6ju6 ^ Hu4ju6));
assign Su6ju6 = (~(Zu6ju6 & Gv6ju6));
assign Gv6ju6 = (Nv6ju6 & Uv6ju6);
assign Uv6ju6 = (~(Kc6ju6 & S8fpw6[5]));
assign Nv6ju6 = (~(S8fpw6[7] & Xv4ju6));
assign Zu6ju6 = (Bw6ju6 & Iw6ju6);
assign Iw6ju6 = (~(Sw4ju6 & Uo6ju6));
assign Bw6ju6 = (Gx4ju6 | Ad8iu6);
assign Nh6ju6 = (~(J1liu6 | Yykiu6));
assign Yykiu6 = (~(Pw6ju6 & Ww6ju6));
assign Ww6ju6 = (Dx6ju6 & Kx6ju6);
assign Kx6ju6 = (~(By4ju6 & Eafpw6[24]));
assign Dx6ju6 = (~(Affpw6[24] | Wk4ju6));
assign Pw6ju6 = (Rx6ju6 & Yx6ju6);
assign Yx6ju6 = (~(Iy4ju6 & Fy6ju6));
assign Rx6ju6 = (Yj0iu6 ? Ty6ju6 : My6ju6);
assign Ty6ju6 = (~(Ys4ju6 & Qbfpw6[24]));
assign My6ju6 = (~(Az6ju6 | Mt4ju6));
assign Az6ju6 = (Qbfpw6[24] ? Tt4ju6 : Ys4ju6);
assign Qbfpw6[24] = (Hz6ju6 | M75ju6);
assign Hz6ju6 = (Fy6ju6 ? A85ju6 : T75ju6);
assign J1liu6 = (~(Oz6ju6 & Vz6ju6));
assign Vz6ju6 = (C07ju6 & J07ju6);
assign J07ju6 = (~(By4ju6 & Eafpw6[26]));
assign C07ju6 = (~(Affpw6[26] | Q07ju6));
assign Q07ju6 = (~(X07ju6 | E17ju6));
assign X07ju6 = (Qbfpw6[26] ? Wc5ju6 : Cg5ju6);
assign Oz6ju6 = (L17ju6 & S17ju6);
assign S17ju6 = (~(Iy4ju6 & Z17ju6));
assign L17ju6 = (~(Ub5ju6 & G27ju6));
assign G27ju6 = (~(N27ju6 & Ic5ju6));
assign N27ju6 = (~(E17ju6 & Qbfpw6[26]));
assign Qbfpw6[26] = (U27ju6 | M75ju6);
assign U27ju6 = (Z17ju6 ? A85ju6 : T75ju6);
assign E17ju6 = (!Kj0iu6);
assign Zg6ju6 = (B37ju6 & I37ju6);
assign I37ju6 = (~(W4liu6 | B4liu6));
assign B4liu6 = (~(P37ju6 & W37ju6));
assign W37ju6 = (D47ju6 & K47ju6);
assign K47ju6 = (~(By4ju6 & Eafpw6[27]));
assign D47ju6 = (~(Affpw6[27] | R47ju6));
assign R47ju6 = (~(Y47ju6 | F57ju6));
assign Y47ju6 = (Qbfpw6[27] ? Wc5ju6 : Cg5ju6);
assign P37ju6 = (M57ju6 & T57ju6);
assign T57ju6 = (~(Iy4ju6 & A67ju6));
assign M57ju6 = (~(Ub5ju6 & H67ju6));
assign H67ju6 = (~(O67ju6 & Ic5ju6));
assign O67ju6 = (~(F57ju6 & Qbfpw6[27]));
assign Qbfpw6[27] = (V67ju6 | M75ju6);
assign V67ju6 = (A67ju6 ? A85ju6 : T75ju6);
assign F57ju6 = (!Dj0iu6);
assign W4liu6 = (~(C77ju6 & J77ju6));
assign J77ju6 = (Q77ju6 & X77ju6);
assign X77ju6 = (~(I55ju6 & vis_apsr_o[1]));
assign Q77ju6 = (~(Affpw6[29] | Wk4ju6));
assign C77ju6 = (E87ju6 & L87ju6);
assign L87ju6 = (Pi0iu6 ? Z87ju6 : S87ju6);
assign Z87ju6 = (~(Ys4ju6 & Qbfpw6[29]));
assign S87ju6 = (~(G97ju6 | Mt4ju6));
assign G97ju6 = (Qbfpw6[29] ? Tt4ju6 : Ys4ju6);
assign Qbfpw6[29] = (N97ju6 | M75ju6);
assign N97ju6 = (Wh8iu6 ? A85ju6 : T75ju6);
assign E87ju6 = (U97ju6 & Ba7ju6);
assign Ba7ju6 = (~(By4ju6 & Eafpw6[29]));
assign U97ju6 = (~(Iy4ju6 & Wh8iu6));
assign B37ju6 = (Kgoiu6 & Bpliu6);
assign Bpliu6 = (Ia7ju6 & Pa7ju6);
assign Pa7ju6 = (Wa7ju6 & Db7ju6);
assign Db7ju6 = (~(Pk4ju6 & vis_ipsr_o[1]));
assign Pk4ju6 = (Kb7ju6 & T05ju6);
assign Kb7ju6 = (~(Je8iu6 | S8fpw6[4]));
assign Wa7ju6 = (~(Affpw6[1] | Rb7ju6));
assign Rb7ju6 = (Yb7ju6 & Fc7ju6);
assign Fc7ju6 = (~(B5kiu6 | Qjoiu6));
assign Yb7ju6 = (vis_control_o & T05ju6);
assign Ia7ju6 = (Mc7ju6 & Tc7ju6);
assign Tc7ju6 = (Hl0iu6 ? Hd7ju6 : Ad7ju6);
assign Hd7ju6 = (~(Ys4ju6 & Qbfpw6[1]));
assign Ad7ju6 = (~(Od7ju6 | Mt4ju6));
assign Od7ju6 = (Qbfpw6[1] ? Tt4ju6 : Ys4ju6);
assign Qbfpw6[1] = (~(Vd7ju6 ^ Hu4ju6));
assign Vd7ju6 = (~(Ce7ju6 & Je7ju6));
assign Je7ju6 = (Rb8iu6 | Gx4ju6);
assign Ce7ju6 = (Qe7ju6 & Xe7ju6);
assign Xe7ju6 = (~(S8fpw6[1] & E35ju6));
assign E35ju6 = (Xv4ju6 | Ef7ju6);
assign Ef7ju6 = (Lf7ju6 & Sf7ju6);
assign Lf7ju6 = (H6ghu6 & Cyfpw6[1]);
assign Xv4ju6 = (Zf7ju6 | Gg7ju6);
assign Gg7ju6 = (H6ghu6 & Ng7ju6);
assign Ng7ju6 = (~(Ug7ju6 & Bh7ju6));
assign Bh7ju6 = (~(Ih7ju6 & K9aiu6));
assign Ih7ju6 = (~(Ph7ju6 & Wh7ju6));
assign Ph7ju6 = (M32ju6 | Cyfpw6[6]);
assign Ug7ju6 = (Di7ju6 & Ki7ju6);
assign Ki7ju6 = (~(Fd0iu6 & Ri7ju6));
assign Ri7ju6 = (Mo2ju6 | Yi7ju6);
assign Di7ju6 = (~(C0ehu6 & Fj7ju6));
assign Fj7ju6 = (~(O60ju6 & Mj7ju6));
assign Mj7ju6 = (~(Jf6ju6 & Cyfpw6[0]));
assign Qe7ju6 = (~(Sw4ju6 & Znliu6));
assign Mc7ju6 = (Tj7ju6 & Ak7ju6);
assign Ak7ju6 = (~(By4ju6 & Eafpw6[1]));
assign Tj7ju6 = (~(Iy4ju6 & Znliu6));
assign Kgoiu6 = (Hk7ju6 & Ok7ju6);
assign Ok7ju6 = (Vk7ju6 & Cl7ju6);
assign Cl7ju6 = (~(vis_apsr_o[0] & I55ju6));
assign I55ju6 = (Jl7ju6 & T05ju6);
assign T05ju6 = (Ql7ju6 & Xl7ju6);
assign Xl7ju6 = (~(Qxaiu6 | C0ehu6));
assign Ql7ju6 = (H6ghu6 & D31ju6);
assign Jl7ju6 = (~(S8fpw6[2] | S8fpw6[4]));
assign Vk7ju6 = (~(Affpw6[28] | Wk4ju6));
assign Hk7ju6 = (Em7ju6 & Lm7ju6);
assign Lm7ju6 = (Wi0iu6 ? Zm7ju6 : Sm7ju6);
assign Zm7ju6 = (~(Ys4ju6 & Qbfpw6[28]));
assign Sm7ju6 = (~(Gn7ju6 | Mt4ju6));
assign Gn7ju6 = (Qbfpw6[28] ? Tt4ju6 : Ys4ju6);
assign Qbfpw6[28] = (Nn7ju6 | M75ju6);
assign Nn7ju6 = (Mbniu6 ? T75ju6 : A85ju6);
assign Em7ju6 = (Un7ju6 & Bo7ju6);
assign Bo7ju6 = (~(By4ju6 & Eafpw6[28]));
assign Un7ju6 = (Io7ju6 | Mbniu6);
assign Mbniu6 = (!Po7ju6);
assign Jh4ju6 = (Wo7ju6 & Dp7ju6);
assign Dp7ju6 = (Kp7ju6 & Rp7ju6);
assign Rp7ju6 = (Yp7ju6 & Fq7ju6);
assign Fq7ju6 = (~(R3niu6 | L7niu6));
assign L7niu6 = (~(Mq7ju6 & Tq7ju6));
assign Tq7ju6 = (Ar7ju6 & Hr7ju6);
assign Hr7ju6 = (~(Or7ju6 & Ub5ju6));
assign Or7ju6 = (~(Ic5ju6 & Vr7ju6));
assign Vr7ju6 = (~(Ve0iu6 & W4epw6));
assign Ar7ju6 = (~(Affpw6[8] | Cs7ju6));
assign Cs7ju6 = (~(Js7ju6 | Ve0iu6));
assign Ve0iu6 = (Mm4ju6 ? Qs7ju6 : Q6niu6);
assign Qs7ju6 = (Xs7ju6 & Et7ju6);
assign Et7ju6 = (Lt7ju6 & St7ju6);
assign St7ju6 = (Zt7ju6 & Gu7ju6);
assign Gu7ju6 = (~(Jo4ju6 & vis_r14_o[8]));
assign Zt7ju6 = (Nu7ju6 & Uu7ju6);
assign Uu7ju6 = (~(Ep4ju6 & vis_psp_o[6]));
assign Nu7ju6 = (~(Lp4ju6 & vis_msp_o[6]));
assign Lt7ju6 = (Bv7ju6 & Iv7ju6);
assign Iv7ju6 = (~(Gq4ju6 & vis_r12_o[8]));
assign Bv7ju6 = (~(Nq4ju6 & vis_r11_o[8]));
assign Xs7ju6 = (Pv7ju6 & Wv7ju6);
assign Wv7ju6 = (Dw7ju6 & Kw7ju6);
assign Kw7ju6 = (~(Wr4ju6 & vis_r10_o[8]));
assign Dw7ju6 = (~(Ds4ju6 & vis_r9_o[8]));
assign Pv7ju6 = (B40iu6 & Rw7ju6);
assign Rw7ju6 = (~(Rs4ju6 & vis_r8_o[8]));
assign Q6niu6 = (!Fkfpw6[8]);
assign Js7ju6 = (W4epw6 ? Wc5ju6 : Cg5ju6);
assign W4epw6 = (~(Yw7ju6 ^ Hu4ju6));
assign Yw7ju6 = (~(Fx7ju6 & Mx7ju6));
assign Mx7ju6 = (Tx7ju6 & Ay7ju6);
assign Ay7ju6 = (~(Kc6ju6 & S8fpw6[6]));
assign Tx7ju6 = (~(Zf7ju6 & S8fpw6[8]));
assign Fx7ju6 = (Hy7ju6 & Oy7ju6);
assign Oy7ju6 = (Vy7ju6 | Cz7ju6);
assign Hy7ju6 = (O95iu6 | Gx4ju6);
assign Mq7ju6 = (Jz7ju6 & Qz7ju6);
assign Qz7ju6 = (~(By4ju6 & Eafpw6[8]));
assign Jz7ju6 = (Io7ju6 | Cz7ju6);
assign R3niu6 = (~(Xz7ju6 & E08ju6));
assign E08ju6 = (L08ju6 & S08ju6);
assign S08ju6 = (~(By4ju6 & Eafpw6[9]));
assign L08ju6 = (~(Affpw6[9] | Z08ju6));
assign Z08ju6 = (~(G18ju6 | N18ju6));
assign G18ju6 = (Q5phu6 ? Wc5ju6 : Cg5ju6);
assign Xz7ju6 = (U18ju6 & B28ju6);
assign B28ju6 = (Io7ju6 | I28ju6);
assign U18ju6 = (~(Ub5ju6 & P28ju6));
assign P28ju6 = (~(W28ju6 & Ic5ju6));
assign W28ju6 = (~(N18ju6 & Q5phu6));
assign Q5phu6 = (D38ju6 ^ Ol6ju6);
assign D38ju6 = (~(K38ju6 & R38ju6));
assign R38ju6 = (Y38ju6 & F48ju6);
assign F48ju6 = (~(Kc6ju6 & S8fpw6[7]));
assign Kc6ju6 = (H6ghu6 & M48ju6);
assign M48ju6 = (~(T48ju6 & A58ju6));
assign A58ju6 = (Cyfpw6[3] ? O58ju6 : H58ju6);
assign O58ju6 = (V58ju6 | Jc2ju6);
assign H58ju6 = (Szniu6 | Knaiu6);
assign T48ju6 = (C68ju6 & J68ju6);
assign J68ju6 = (~(Y2aiu6 & Vo3ju6));
assign Y2aiu6 = (Q68ju6 & Fd0iu6);
assign Q68ju6 = (~(As0iu6 | C0ehu6));
assign C68ju6 = (~(D6kiu6 & X68ju6));
assign X68ju6 = (~(E78ju6 & Jc2ju6));
assign E78ju6 = (~(L78ju6 | Cyfpw6[3]));
assign Y38ju6 = (~(Zf7ju6 & S8fpw6[9]));
assign K38ju6 = (S78ju6 & Z78ju6);
assign Z78ju6 = (Vy7ju6 | I28ju6);
assign S78ju6 = (Ndiiu6 | Gx4ju6);
assign N18ju6 = (!He0iu6);
assign Yp7ju6 = (~(Vsliu6 | Vymiu6));
assign Vymiu6 = (~(G88ju6 & N88ju6));
assign N88ju6 = (U88ju6 & B98ju6);
assign B98ju6 = (~(By4ju6 & Eafpw6[10]));
assign U88ju6 = (~(Affpw6[10] | I98ju6));
assign I98ju6 = (~(P98ju6 | Zn0iu6));
assign P98ju6 = (Qbfpw6[10] ? Wc5ju6 : Cg5ju6);
assign G88ju6 = (W98ju6 & Da8ju6);
assign Da8ju6 = (Io7ju6 | Ka8ju6);
assign Io7ju6 = (!Iy4ju6);
assign W98ju6 = (~(Ub5ju6 & Ra8ju6));
assign Ra8ju6 = (~(Ya8ju6 & Ic5ju6));
assign Ya8ju6 = (~(Zn0iu6 & Qbfpw6[10]));
assign Qbfpw6[10] = (~(Fb8ju6 ^ Hu4ju6));
assign Fb8ju6 = (~(Mb8ju6 & Tb8ju6));
assign Tb8ju6 = (Tniiu6 | Gx4ju6);
assign Mb8ju6 = (Ac8ju6 & Hc8ju6);
assign Hc8ju6 = (~(Zf7ju6 & S8fpw6[10]));
assign Ac8ju6 = (Vy7ju6 | Ka8ju6);
assign Zn0iu6 = (Cn5ju6 ? Aymiu6 : Oc8ju6);
assign Aymiu6 = (!Fkfpw6[10]);
assign Oc8ju6 = (Vc8ju6 & Cd8ju6);
assign Cd8ju6 = (Jd8ju6 & Qd8ju6);
assign Qd8ju6 = (Xd8ju6 & Ee8ju6);
assign Ee8ju6 = (~(Jo4ju6 & vis_r14_o[10]));
assign Xd8ju6 = (Le8ju6 & Se8ju6);
assign Se8ju6 = (~(Ep4ju6 & vis_psp_o[8]));
assign Le8ju6 = (~(Lp4ju6 & vis_msp_o[8]));
assign Jd8ju6 = (Ze8ju6 & Gf8ju6);
assign Gf8ju6 = (~(Gq4ju6 & vis_r12_o[10]));
assign Ze8ju6 = (~(Nq4ju6 & vis_r11_o[10]));
assign Vc8ju6 = (Nf8ju6 & Uf8ju6);
assign Uf8ju6 = (Bg8ju6 & Ig8ju6);
assign Ig8ju6 = (~(Wr4ju6 & vis_r10_o[10]));
assign Bg8ju6 = (~(Ds4ju6 & vis_r9_o[10]));
assign Nf8ju6 = (Wb0iu6 & Pg8ju6);
assign Pg8ju6 = (~(Rs4ju6 & vis_r8_o[10]));
assign Vsliu6 = (~(Wg8ju6 & Dh8ju6));
assign Dh8ju6 = (Kh8ju6 & Rh8ju6);
assign Rh8ju6 = (~(By4ju6 & Eafpw6[25]));
assign Kh8ju6 = (~(Affpw6[25] | Yh8ju6));
assign Yh8ju6 = (~(Fi8ju6 | Mi8ju6));
assign Fi8ju6 = (Qbfpw6[25] ? Wc5ju6 : Cg5ju6);
assign Wg8ju6 = (Ti8ju6 & Aj8ju6);
assign Aj8ju6 = (~(Iy4ju6 & Goliu6));
assign Ti8ju6 = (~(Ub5ju6 & Hj8ju6));
assign Hj8ju6 = (~(Oj8ju6 & Ic5ju6));
assign Oj8ju6 = (~(Mi8ju6 & Qbfpw6[25]));
assign Qbfpw6[25] = (Vj8ju6 | M75ju6);
assign M75ju6 = (~(Ck8ju6 & Jk8ju6));
assign Jk8ju6 = (~(T75ju6 & Vy7ju6));
assign Ck8ju6 = (~(Hu4ju6 & Qk8ju6));
assign Qk8ju6 = (~(Xk8ju6 & Ij5ju6));
assign Vj8ju6 = (Goliu6 ? A85ju6 : T75ju6);
assign A85ju6 = (~(Vy7ju6 | Ol6ju6));
assign T75ju6 = (El8ju6 & Ol6ju6);
assign Ol6ju6 = (!Hu4ju6);
assign El8ju6 = (Xk8ju6 & Ij5ju6);
assign Mi8ju6 = (!Rj0iu6);
assign Kp7ju6 = (Ll8ju6 & Sl8ju6);
assign Sl8ju6 = (~(Pomiu6 | Bvmiu6));
assign Bvmiu6 = (~(Zl8ju6 & Gm8ju6));
assign Gm8ju6 = (Nm8ju6 & Um8ju6);
assign Um8ju6 = (~(By4ju6 & Eafpw6[11]));
assign Nm8ju6 = (~(Affpw6[11] | Bn8ju6));
assign Bn8ju6 = (Iy4ju6 & In8ju6);
assign Zl8ju6 = (Pn8ju6 & Wn8ju6);
assign Wn8ju6 = (~(Ub5ju6 & Do8ju6));
assign Do8ju6 = (~(Ko8ju6 & Ic5ju6));
assign Ko8ju6 = (~(Sn0iu6 & C1epw6));
assign Pn8ju6 = (Ro8ju6 | Sn0iu6);
assign Sn0iu6 = (Cn5ju6 ? Ormiu6 : Yo8ju6);
assign Ormiu6 = (!Fkfpw6[11]);
assign Yo8ju6 = (Fp8ju6 & Mp8ju6);
assign Mp8ju6 = (Tp8ju6 & Aq8ju6);
assign Aq8ju6 = (Hq8ju6 & Oq8ju6);
assign Oq8ju6 = (~(Jo4ju6 & vis_r14_o[11]));
assign Hq8ju6 = (Vq8ju6 & Cr8ju6);
assign Cr8ju6 = (~(Ep4ju6 & vis_psp_o[9]));
assign Vq8ju6 = (~(Lp4ju6 & vis_msp_o[9]));
assign Tp8ju6 = (Jr8ju6 & Qr8ju6);
assign Qr8ju6 = (~(Gq4ju6 & vis_r12_o[11]));
assign Jr8ju6 = (~(Nq4ju6 & vis_r11_o[11]));
assign Fp8ju6 = (Xr8ju6 & Es8ju6);
assign Es8ju6 = (Ls8ju6 & Ss8ju6);
assign Ss8ju6 = (~(Wr4ju6 & vis_r10_o[11]));
assign Ls8ju6 = (~(Ds4ju6 & vis_r9_o[11]));
assign Xr8ju6 = (Pb0iu6 & Zs8ju6);
assign Zs8ju6 = (~(Rs4ju6 & vis_r8_o[11]));
assign Ro8ju6 = (C1epw6 ? Wc5ju6 : Cg5ju6);
assign C1epw6 = (~(Gt8ju6 ^ Hu4ju6));
assign Gt8ju6 = (~(Nt8ju6 & Ut8ju6));
assign Ut8ju6 = (I6jiu6 | Gx4ju6);
assign Nt8ju6 = (Bu8ju6 & Ij5ju6);
assign Bu8ju6 = (~(Sw4ju6 & In8ju6));
assign Pomiu6 = (~(Iu8ju6 & Pu8ju6));
assign Pu8ju6 = (Wu8ju6 & Dv8ju6);
assign Dv8ju6 = (~(By4ju6 & Eafpw6[12]));
assign Wu8ju6 = (~(Affpw6[12] | Kv8ju6));
assign Kv8ju6 = (Iy4ju6 & Rv8ju6);
assign Iu8ju6 = (Yv8ju6 & Fw8ju6);
assign Fw8ju6 = (~(Ub5ju6 & Mw8ju6));
assign Mw8ju6 = (~(Tw8ju6 & Ic5ju6));
assign Tw8ju6 = (~(Ln0iu6 & J1epw6));
assign Yv8ju6 = (Ax8ju6 | Ln0iu6);
assign Ax8ju6 = (J1epw6 ? Wc5ju6 : Cg5ju6);
assign J1epw6 = (~(Hx8ju6 ^ Hu4ju6));
assign Hx8ju6 = (~(Ox8ju6 & Vx8ju6));
assign Vx8ju6 = (Y8biu6 | Gx4ju6);
assign Ox8ju6 = (Cy8ju6 & Ij5ju6);
assign Cy8ju6 = (~(Sw4ju6 & Rv8ju6));
assign Ll8ju6 = (~(Fjmiu6 | Xlmiu6));
assign Xlmiu6 = (~(Jy8ju6 & Qy8ju6));
assign Qy8ju6 = (Xy8ju6 & Ez8ju6);
assign Ez8ju6 = (~(By4ju6 & Eafpw6[13]));
assign Xy8ju6 = (~(Affpw6[13] | Lz8ju6));
assign Lz8ju6 = (Iy4ju6 & Sz8ju6);
assign Jy8ju6 = (Zz8ju6 & G09ju6);
assign G09ju6 = (~(Ub5ju6 & N09ju6));
assign N09ju6 = (~(U09ju6 & Ic5ju6));
assign U09ju6 = (~(En0iu6 & Q1epw6));
assign Zz8ju6 = (B19ju6 | En0iu6);
assign B19ju6 = (Q1epw6 ? Wc5ju6 : Cg5ju6);
assign Q1epw6 = (~(I19ju6 ^ Hu4ju6));
assign I19ju6 = (~(P19ju6 & W19ju6));
assign W19ju6 = (B5kiu6 | Gx4ju6);
assign P19ju6 = (D29ju6 & Ij5ju6);
assign D29ju6 = (~(Sw4ju6 & Sz8ju6));
assign Fjmiu6 = (~(K29ju6 & R29ju6));
assign R29ju6 = (Y29ju6 & F39ju6);
assign F39ju6 = (~(By4ju6 & Eafpw6[14]));
assign Y29ju6 = (~(Affpw6[14] | M39ju6));
assign M39ju6 = (Iy4ju6 & T39ju6);
assign K29ju6 = (A49ju6 & H49ju6);
assign H49ju6 = (~(Ub5ju6 & O49ju6));
assign O49ju6 = (~(V49ju6 & Ic5ju6));
assign V49ju6 = (~(Xm0iu6 & X1epw6));
assign A49ju6 = (C59ju6 | Xm0iu6);
assign C59ju6 = (X1epw6 ? Wc5ju6 : Cg5ju6);
assign X1epw6 = (~(J59ju6 ^ Hu4ju6));
assign J59ju6 = (~(Q59ju6 & X59ju6));
assign X59ju6 = (Gx4ju6 | Cajiu6);
assign Q59ju6 = (E69ju6 & Ij5ju6);
assign E69ju6 = (~(Sw4ju6 & T39ju6));
assign Wo7ju6 = (L69ju6 & S69ju6);
assign S69ju6 = (Z69ju6 & G79ju6);
assign G79ju6 = (Vdmiu6 & Ngmiu6);
assign Ngmiu6 = (N79ju6 & U79ju6);
assign U79ju6 = (B89ju6 & I89ju6);
assign I89ju6 = (~(By4ju6 & Eafpw6[15]));
assign B89ju6 = (~(Affpw6[15] | P89ju6));
assign P89ju6 = (Iy4ju6 & W89ju6);
assign N79ju6 = (D99ju6 & K99ju6);
assign K99ju6 = (~(Ub5ju6 & R99ju6));
assign R99ju6 = (~(Y99ju6 & Ic5ju6));
assign Y99ju6 = (~(Qm0iu6 & L2epw6));
assign D99ju6 = (Fa9ju6 | Qm0iu6);
assign Fa9ju6 = (L2epw6 ? Wc5ju6 : Cg5ju6);
assign L2epw6 = (~(Ma9ju6 ^ Hu4ju6));
assign Ma9ju6 = (~(Ta9ju6 & Ab9ju6));
assign Ab9ju6 = (Gx4ju6 | Qjoiu6);
assign Ta9ju6 = (Hb9ju6 & Ij5ju6);
assign Hb9ju6 = (~(Sw4ju6 & W89ju6));
assign Vdmiu6 = (Ob9ju6 & Vb9ju6);
assign Vb9ju6 = (Cc9ju6 & Jc9ju6);
assign Jc9ju6 = (~(By4ju6 & Eafpw6[16]));
assign Cc9ju6 = (~(Affpw6[16] | Qc9ju6));
assign Qc9ju6 = (Iy4ju6 & Xc9ju6);
assign Ob9ju6 = (Ed9ju6 & Ld9ju6);
assign Ld9ju6 = (~(Ub5ju6 & Sd9ju6));
assign Sd9ju6 = (~(Zd9ju6 & Ic5ju6));
assign Zd9ju6 = (~(Jm0iu6 & Z2epw6));
assign Ed9ju6 = (Ge9ju6 | Jm0iu6);
assign Ge9ju6 = (Z2epw6 ? Wc5ju6 : Cg5ju6);
assign Z2epw6 = (~(Ne9ju6 ^ Hu4ju6));
assign Ne9ju6 = (~(Ue9ju6 & Bf9ju6));
assign Bf9ju6 = (~(If9ju6 & S8fpw6[5]));
assign Ue9ju6 = (Pf9ju6 & Ij5ju6);
assign Pf9ju6 = (~(Sw4ju6 & Xc9ju6));
assign Z69ju6 = (X7miu6 & Wamiu6);
assign Wamiu6 = (Wf9ju6 & Dg9ju6);
assign Dg9ju6 = (Kg9ju6 & Rg9ju6);
assign Rg9ju6 = (~(By4ju6 & Eafpw6[17]));
assign Kg9ju6 = (~(Affpw6[17] | Yg9ju6));
assign Yg9ju6 = (Iy4ju6 & Fh9ju6);
assign Wf9ju6 = (Mh9ju6 & Th9ju6);
assign Th9ju6 = (~(Ub5ju6 & Ai9ju6));
assign Ai9ju6 = (~(Hi9ju6 & Ic5ju6));
assign Hi9ju6 = (~(Cm0iu6 & G3epw6));
assign Mh9ju6 = (Oi9ju6 | Cm0iu6);
assign Oi9ju6 = (G3epw6 ? Wc5ju6 : Cg5ju6);
assign G3epw6 = (~(Vi9ju6 ^ Hu4ju6));
assign Vi9ju6 = (~(Cj9ju6 & Jj9ju6));
assign Jj9ju6 = (~(If9ju6 & S8fpw6[6]));
assign Cj9ju6 = (Qj9ju6 & Ij5ju6);
assign Qj9ju6 = (~(Sw4ju6 & Fh9ju6));
assign X7miu6 = (Xj9ju6 & Ek9ju6);
assign Ek9ju6 = (Lk9ju6 & Sk9ju6);
assign Sk9ju6 = (~(By4ju6 & Eafpw6[18]));
assign Lk9ju6 = (~(Affpw6[18] | Zk9ju6));
assign Zk9ju6 = (Iy4ju6 & Gl9ju6);
assign Xj9ju6 = (Nl9ju6 & Ul9ju6);
assign Ul9ju6 = (~(Ub5ju6 & Bm9ju6));
assign Bm9ju6 = (~(Im9ju6 & Ic5ju6));
assign Im9ju6 = (~(Vl0iu6 & N3epw6));
assign Nl9ju6 = (Pm9ju6 | Vl0iu6);
assign Pm9ju6 = (N3epw6 ? Wc5ju6 : Cg5ju6);
assign N3epw6 = (~(Wm9ju6 ^ Hu4ju6));
assign Wm9ju6 = (~(Dn9ju6 & Kn9ju6));
assign Kn9ju6 = (~(If9ju6 & S8fpw6[7]));
assign Dn9ju6 = (Rn9ju6 & Ij5ju6);
assign Rn9ju6 = (~(Sw4ju6 & Gl9ju6));
assign L69ju6 = (Yn9ju6 & Fo9ju6);
assign Fo9ju6 = (Z1miu6 & Y4miu6);
assign Y4miu6 = (Mo9ju6 & To9ju6);
assign To9ju6 = (Ap9ju6 & Hp9ju6);
assign Hp9ju6 = (~(By4ju6 & Eafpw6[19]));
assign Ap9ju6 = (~(Affpw6[19] | Op9ju6));
assign Op9ju6 = (Iy4ju6 & Vp9ju6);
assign Mo9ju6 = (Cq9ju6 & Jq9ju6);
assign Jq9ju6 = (~(Ub5ju6 & Qq9ju6));
assign Qq9ju6 = (~(Xq9ju6 & Ic5ju6));
assign Xq9ju6 = (~(Ol0iu6 & U3epw6));
assign Cq9ju6 = (Er9ju6 | Ol0iu6);
assign Er9ju6 = (U3epw6 ? Wc5ju6 : Cg5ju6);
assign U3epw6 = (~(Lr9ju6 ^ Hu4ju6));
assign Lr9ju6 = (~(Sr9ju6 & Zr9ju6));
assign Zr9ju6 = (Gx4ju6 | I65iu6);
assign Sr9ju6 = (Gs9ju6 & Ij5ju6);
assign Gs9ju6 = (~(Sw4ju6 & Vp9ju6));
assign Z1miu6 = (Ns9ju6 & Us9ju6);
assign Us9ju6 = (Bt9ju6 & It9ju6);
assign It9ju6 = (~(By4ju6 & Eafpw6[20]));
assign Bt9ju6 = (~(Affpw6[20] | Pt9ju6));
assign Pt9ju6 = (Iy4ju6 & Wt9ju6);
assign Ns9ju6 = (Du9ju6 & Ku9ju6);
assign Ku9ju6 = (~(Ub5ju6 & Ru9ju6));
assign Ru9ju6 = (~(Yu9ju6 & Ic5ju6));
assign Yu9ju6 = (~(Al0iu6 & B4epw6));
assign Du9ju6 = (Fv9ju6 | Al0iu6);
assign Fv9ju6 = (B4epw6 ? Wc5ju6 : Cg5ju6);
assign B4epw6 = (~(Mv9ju6 ^ Hu4ju6));
assign Mv9ju6 = (~(Tv9ju6 & Aw9ju6));
assign Aw9ju6 = (Gx4ju6 | P65iu6);
assign Tv9ju6 = (Hw9ju6 & Ij5ju6);
assign Hw9ju6 = (~(Sw4ju6 & Wt9ju6));
assign Yn9ju6 = (Uvliu6 & Azliu6);
assign Azliu6 = (Ow9ju6 & Vw9ju6);
assign Vw9ju6 = (Cx9ju6 & Jx9ju6);
assign Jx9ju6 = (~(By4ju6 & Eafpw6[21]));
assign Cx9ju6 = (~(Affpw6[21] | Qx9ju6));
assign Qx9ju6 = (Iy4ju6 & Xx9ju6);
assign Ow9ju6 = (Ey9ju6 & Ly9ju6);
assign Ly9ju6 = (~(Ub5ju6 & Sy9ju6));
assign Sy9ju6 = (~(Zy9ju6 & Ic5ju6));
assign Zy9ju6 = (~(Tk0iu6 & I4epw6));
assign Ey9ju6 = (Gz9ju6 | Tk0iu6);
assign Gz9ju6 = (I4epw6 ? Wc5ju6 : Cg5ju6);
assign I4epw6 = (~(Nz9ju6 ^ Hu4ju6));
assign Nz9ju6 = (~(Uz9ju6 & B0aju6));
assign B0aju6 = (~(If9ju6 & S8fpw6[10]));
assign Uz9ju6 = (I0aju6 & Ij5ju6);
assign I0aju6 = (~(Sw4ju6 & Xx9ju6));
assign Uvliu6 = (P0aju6 & W0aju6);
assign W0aju6 = (D1aju6 & K1aju6);
assign K1aju6 = (~(By4ju6 & Eafpw6[22]));
assign By4ju6 = (H6ghu6 & R1aju6);
assign R1aju6 = (Y1aju6 | Pt2ju6);
assign Y1aju6 = (Cyfpw6[4] ? Difiu6 : F2aju6);
assign F2aju6 = (~(M2aju6 & T2aju6));
assign T2aju6 = (Qcoiu6 | H4ghu6);
assign M2aju6 = (~(A3aju6 | H3aju6));
assign D1aju6 = (~(Affpw6[22] | O3aju6));
assign O3aju6 = (Iy4ju6 & V3aju6);
assign Iy4ju6 = (H6ghu6 & C4aju6);
assign C4aju6 = (J4aju6 | S6aiu6);
assign P0aju6 = (Q4aju6 & X4aju6);
assign X4aju6 = (~(Ub5ju6 & E5aju6));
assign E5aju6 = (~(L5aju6 & Ic5ju6));
assign L5aju6 = (~(Mk0iu6 & P4epw6));
assign Ub5ju6 = (Wk4ju6 | Ys4ju6);
assign Wk4ju6 = (!Ic5ju6);
assign Ic5ju6 = (~(S5aju6 & H6ghu6));
assign S5aju6 = (Md0iu6 & H4ghu6);
assign Q4aju6 = (Z5aju6 | Mk0iu6);
assign Z5aju6 = (P4epw6 ? Wc5ju6 : Cg5ju6);
assign P4epw6 = (~(G6aju6 ^ Hu4ju6));
assign Hu4ju6 = (~(H6ghu6 & N6aju6));
assign N6aju6 = (~(U6aju6 & B7aju6));
assign B7aju6 = (I7aju6 & P7aju6);
assign P7aju6 = (~(W7aju6 & Cyfpw6[4]));
assign W7aju6 = (D8aju6 & Hs0iu6);
assign D8aju6 = (~(Wfoiu6 & K8aju6));
assign K8aju6 = (Tr0iu6 | Cyfpw6[6]);
assign I7aju6 = (R8aju6 & Zu0iu6);
assign Zu0iu6 = (~(Y8aju6 & F9aju6));
assign R8aju6 = (~(M9aju6 & A3aju6));
assign M9aju6 = (S2ziu6 & C0ehu6);
assign U6aju6 = (Lu0iu6 & T9aju6);
assign T9aju6 = (~(Bi0iu6 & Tfjiu6));
assign Lu0iu6 = (Aaaju6 & Haaju6);
assign Haaju6 = (Ey2ju6 | Ezniu6);
assign Ezniu6 = (!F23ju6);
assign Aaaju6 = (Oaaju6 & Vaaju6);
assign Vaaju6 = (~(Mo2ju6 & C0ehu6));
assign Oaaju6 = (~(L78ju6 & D6kiu6));
assign G6aju6 = (~(Cbaju6 & Jbaju6));
assign Jbaju6 = (D7fpw6[11] ? Xk8ju6 : Qbaju6);
assign Xk8ju6 = (!Ui5ju6);
assign Ui5ju6 = (If9ju6 & S8fpw6[11]);
assign Qbaju6 = (Gx4ju6 | S8fpw6[11]);
assign Gx4ju6 = (!If9ju6);
assign If9ju6 = (Xbaju6 & Sy2ju6);
assign Xbaju6 = (H6ghu6 & Fd0iu6);
assign Cbaju6 = (Ecaju6 & Ij5ju6);
assign Ij5ju6 = (~(Zf7ju6 & S8fpw6[11]));
assign Zf7ju6 = (Lcaju6 & H6ghu6);
assign Lcaju6 = (Pt2ju6 & Hzziu6);
assign Ecaju6 = (~(Sw4ju6 & V3aju6));
assign Sw4ju6 = (!Vy7ju6);
assign Vy7ju6 = (~(H6ghu6 & Scaju6));
assign Scaju6 = (~(Zcaju6 & Gdaju6));
assign Gdaju6 = (Ndaju6 & Udaju6);
assign Udaju6 = (~(H4ghu6 & Beaju6));
assign Beaju6 = (~(Ieaju6 & Peaju6));
assign Peaju6 = (~(Owoiu6 | Kfiiu6));
assign Ieaju6 = (Weaju6 & Dfaju6);
assign Dfaju6 = (Wfoiu6 | Vwaiu6);
assign Weaju6 = (Y2oiu6 | Ii0iu6);
assign Ndaju6 = (Kfaju6 & Rfaju6);
assign Rfaju6 = (~(Yfaju6 & Whfiu6));
assign Yfaju6 = (Oiaiu6 & Sq3ju6);
assign Kfaju6 = (~(Cyfpw6[3] & Fgaju6));
assign Fgaju6 = (~(Yn2ju6 & Mgaju6));
assign Mgaju6 = (Z6oiu6 | Wfoiu6);
assign Zcaju6 = (Tgaju6 & Ahaju6);
assign Ahaju6 = (~(Pt2ju6 & Pthiu6));
assign Tgaju6 = (Y2oiu6 | Cyfpw6[7]);
assign Wc5ju6 = (~(Tt4ju6 | Mt4ju6));
assign Tt4ju6 = (~(Hhaju6 & Ohaju6));
assign Ohaju6 = (~(Vhaju6 & H4ghu6));
assign Vhaju6 = (Ciaju6 & Tr0iu6);
assign Ciaju6 = (Hs0iu6 | Kfiiu6);
assign Hhaju6 = (Szniu6 | Wfoiu6);
assign Cg5ju6 = (~(Ys4ju6 | Mt4ju6));
assign Mt4ju6 = (H6ghu6 & Jiaju6);
assign Jiaju6 = (~(Qiaju6 & Xiaju6));
assign Qiaju6 = (Ejaju6 & Ljaju6);
assign Ljaju6 = (~(Ae0iu6 & N3ziu6));
assign Ejaju6 = (Cyfpw6[6] ? Zjaju6 : Sjaju6);
assign Zjaju6 = (Y2oiu6 | R75iu6);
assign Sjaju6 = (Yn2ju6 | Cyfpw6[4]);
assign Ys4ju6 = (Gkaju6 & Nkaju6);
assign Nkaju6 = (~(Y2oiu6 | Cyfpw6[7]));
assign Gkaju6 = (H6ghu6 & Qyniu6);
assign Xe0ju6 = (!Nzoiu6);
assign Nzoiu6 = (I6jiu6 & Oviiu6);
assign Utohu6 = (!Ukaju6);
assign Ukaju6 = (HREADY ? Blaju6 : Ii0iu6);
assign Blaju6 = (Ilaju6 & Plaju6);
assign Plaju6 = (Wlaju6 & Dmaju6);
assign Dmaju6 = (Kmaju6 & Rmaju6);
assign Rmaju6 = (~(Ymaju6 & Eoyiu6));
assign Ymaju6 = (~(H3piu6 | Lkaiu6));
assign Kmaju6 = (Fnaju6 & Mnaju6);
assign Mnaju6 = (~(Tnaju6 & W8aiu6));
assign Tnaju6 = (Cyfpw6[3] & Aoaju6);
assign Aoaju6 = (~(Hoaju6 & Ooaju6));
assign Ooaju6 = (Voaju6 & T0hhu6);
assign Voaju6 = (~(Ftjiu6 | D7fpw6[3]));
assign Hoaju6 = (~(Rg2ju6 | Q5aiu6));
assign Fnaju6 = (~(Cpaju6 & Jpaju6));
assign Jpaju6 = (~(Qpaju6 | D7fpw6[10]));
assign Cpaju6 = (D7fpw6[8] & J9kiu6);
assign Wlaju6 = (Xpaju6 & Eqaju6);
assign Eqaju6 = (~(Wwziu6 & Lqaju6));
assign Lqaju6 = (~(Y2oiu6 & Sqaju6));
assign Sqaju6 = (Zqaju6 | Cyfpw6[5]);
assign Xpaju6 = (Graju6 & Nraju6);
assign Nraju6 = (~(Btoiu6 & Uraju6));
assign Uraju6 = (~(Ctziu6 & Bsaju6));
assign Bsaju6 = (~(U98iu6 & Xe8iu6));
assign Btoiu6 = (~(Cyfpw6[1] | H4ghu6));
assign Graju6 = (~(Isaju6 & F23ju6));
assign Isaju6 = (Frziu6 & Qe8iu6);
assign Ilaju6 = (Psaju6 & Wsaju6);
assign Wsaju6 = (Dtaju6 & K76ow6);
assign K76ow6 = (P5kiu6 | Sijiu6);
assign Dtaju6 = (R76ow6 & Y76ow6);
assign Y76ow6 = (Ctziu6 | V58ju6);
assign V58ju6 = (!F86ow6);
assign Ctziu6 = (Jcaiu6 | R75iu6);
assign R76ow6 = (~(M86ow6 & Tfjiu6));
assign M86ow6 = (~(T86ow6 & A96ow6));
assign A96ow6 = (~(H96ow6 & W8aiu6));
assign H96ow6 = (~(O96ow6 | Cyfpw6[5]));
assign T86ow6 = (V96ow6 & P5kiu6);
assign P5kiu6 = (!Lijiu6);
assign Lijiu6 = (Whfiu6 & Y7ghu6);
assign V96ow6 = (~(Ca6ow6 & Ae0iu6));
assign Ca6ow6 = (U4kiu6 & I30ju6);
assign Psaju6 = (Ja6ow6 & Qa6ow6);
assign Qa6ow6 = (Xa6ow6 | Jcaiu6);
assign Ja6ow6 = (~(Eb6ow6 & Zraiu6));
assign Eb6ow6 = (~(Lb6ow6 & Sb6ow6));
assign Sb6ow6 = (Zb6ow6 & Gc6ow6);
assign Gc6ow6 = (Nc6ow6 & Kb0ju6);
assign Kb0ju6 = (~(Nyiiu6 & Mtjiu6));
assign Nc6ow6 = (Xs0ju6 & Xl0ju6);
assign Zb6ow6 = (Uc6ow6 & Bd6ow6);
assign Bd6ow6 = (~(Dxziu6 & Id6ow6));
assign Id6ow6 = (~(Pd6ow6 & Wd6ow6));
assign Wd6ow6 = (~(De6ow6 & Frziu6));
assign Uc6ow6 = (Ke6ow6 & Re6ow6);
assign Ke6ow6 = (~(Ye6ow6 & Cyfpw6[0]));
assign Ye6ow6 = (Omyiu6 & Ff6ow6);
assign Ff6ow6 = (Tr0iu6 | D31ju6);
assign Lb6ow6 = (Mf6ow6 & Tf6ow6);
assign Tf6ow6 = (Ag6ow6 & Hg6ow6);
assign Hg6ow6 = (~(Il3ju6 & A95iu6));
assign Ag6ow6 = (Og6ow6 & Vg6ow6);
assign Vg6ow6 = (~(Evyiu6 & D7fpw6[15]));
assign Og6ow6 = (~(N3ziu6 & Xzmiu6));
assign Mf6ow6 = (Ch6ow6 & Jh6ow6);
assign Jh6ow6 = (C0ehu6 ? Xh6ow6 : Qh6ow6);
assign Xh6ow6 = (Ei6ow6 & Li6ow6);
assign Li6ow6 = (Si6ow6 & Zi6ow6);
assign Zi6ow6 = (Gj6ow6 & Geaiu6);
assign Gj6ow6 = (Nj6ow6 | D7fpw6[11]);
assign Si6ow6 = (Uj6ow6 & Bk6ow6);
assign Bk6ow6 = (~(Ik6ow6 & D7fpw6[9]));
assign Ik6ow6 = (D7fpw6[7] ? Wk6ow6 : Pk6ow6);
assign Wk6ow6 = (~(Dl6ow6 & Kl6ow6));
assign Kl6ow6 = (~(Y40ju6 & D7fpw6[6]));
assign Dl6ow6 = (Oviiu6 | Gaziu6);
assign Pk6ow6 = (~(Gkiiu6 | D7fpw6[6]));
assign Uj6ow6 = (~(Rl6ow6 & Ftjiu6));
assign Rl6ow6 = (Yl6ow6 | Fm6ow6);
assign Fm6ow6 = (~(O7ziu6 | X1ziu6));
assign Yl6ow6 = (D7fpw6[13] ? D7fpw6[12] : Mm6ow6);
assign Mm6ow6 = (~(Tm6ow6 & An6ow6));
assign Tm6ow6 = (~(X8ziu6 | Jwiiu6));
assign Ei6ow6 = (Hn6ow6 & Y31ju6);
assign Hn6ow6 = (On6ow6 & Vn6ow6);
assign Vn6ow6 = (Co6ow6 | Xuyiu6);
assign Xuyiu6 = (~(Jo6ow6 | Qo6ow6));
assign Qo6ow6 = (D7fpw6[5] ? Xo6ow6 : Kcziu6);
assign Xo6ow6 = (O95iu6 | Ad8iu6);
assign Jo6ow6 = (~(D7fpw6[8] & D7fpw6[9]));
assign On6ow6 = (~(Qxoiu6 & D7fpw6[12]));
assign Qh6ow6 = (~(Ep6ow6 & F23ju6));
assign Ch6ow6 = (Lp6ow6 & Sp6ow6);
assign Sp6ow6 = (~(Pthiu6 & S6aiu6));
assign Lp6ow6 = (H95iu6 | D7fpw6[11]);
assign Ntohu6 = (G81ju6 ? H2fpw6[0] : Zp6ow6);
assign Zp6ow6 = (~(Gq6ow6 & Nq6ow6));
assign Nq6ow6 = (Uq6ow6 & Br6ow6);
assign Br6ow6 = (~(Fb1ju6 & D7fpw6[8]));
assign Uq6ow6 = (~(P91ju6 & D7fpw6[3]));
assign Gq6ow6 = (Ir6ow6 & Pr6ow6);
assign Pr6ow6 = (~(D7fpw6[0] & Ac1ju6));
assign Gtohu6 = (~(Wr6ow6 & Ds6ow6));
assign Ds6ow6 = (Ks6ow6 & Rs6ow6);
assign Rs6ow6 = (~(Egziu6 & Eafpw6[1]));
assign Ks6ow6 = (Ys6ow6 & Sgziu6);
assign Ys6ow6 = (Ft6ow6 | Njciu6);
assign Njciu6 = (Mt6ow6 & Tt6ow6);
assign Tt6ow6 = (Au6ow6 & Hu6ow6);
assign Hu6ow6 = (Cfliu6 | Ou6ow6);
assign Au6ow6 = (Vu6ow6 & Mdliu6);
assign Vu6ow6 = (~(Qfliu6 & Cv6ow6));
assign Mt6ow6 = (Jv6ow6 & Qv6ow6);
assign Qv6ow6 = (Ycliu6 | Xv6ow6);
assign Jv6ow6 = (~(Aeliu6 & Ew6ow6));
assign Wr6ow6 = (Lw6ow6 & Sw6ow6);
assign Sw6ow6 = (~(Zsfpw6[0] & Cmziu6));
assign Lw6ow6 = (Zkhiu6 | Ar8iu6);
assign Zkhiu6 = (!vis_pc_o[0]);
assign Zsohu6 = (!Zw6ow6);
assign Zw6ow6 = (HREADY ? Gx6ow6 : Mr0iu6);
assign Gx6ow6 = (Nx6ow6 & Ux6ow6);
assign Ux6ow6 = (By6ow6 & Iy6ow6);
assign Iy6ow6 = (Py6ow6 & Wy6ow6);
assign Wy6ow6 = (Dz6ow6 & X5aiu6);
assign Py6ow6 = (Kz6ow6 & Rz6ow6);
assign By6ow6 = (Yz6ow6 & F07ow6);
assign F07ow6 = (B1aiu6 & Uloiu6);
assign Yz6ow6 = (M07ow6 & T07ow6);
assign T07ow6 = (~(A17ow6 & Cyfpw6[4]));
assign A17ow6 = (Cyfpw6[5] & H17ow6);
assign H17ow6 = (~(R2aiu6 & O17ow6));
assign O17ow6 = (~(Ae0iu6 & D6kiu6));
assign M07ow6 = (~(V17ow6 & Htyiu6));
assign V17ow6 = (~(C27ow6 | D7fpw6[14]));
assign Nx6ow6 = (J27ow6 & Q27ow6);
assign Q27ow6 = (X27ow6 & E37ow6);
assign E37ow6 = (L37ow6 & S37ow6);
assign S37ow6 = (~(Z37ow6 & K2aiu6));
assign Z37ow6 = (~(Sijiu6 | Kq0iu6));
assign L37ow6 = (Jojiu6 | E62ju6);
assign E62ju6 = (!G47ow6);
assign X27ow6 = (N47ow6 & U47ow6);
assign U47ow6 = (~(B57ow6 & Ii0iu6));
assign B57ow6 = (~(I57ow6 & P57ow6));
assign P57ow6 = (Yn2ju6 | K9aiu6);
assign I57ow6 = (W57ow6 & D67ow6);
assign D67ow6 = (~(K67ow6 & Ae0iu6));
assign K67ow6 = (I30ju6 & Y2oiu6);
assign W57ow6 = (E45iu6 | L62ju6);
assign N47ow6 = (~(R67ow6 & Geaiu6));
assign R67ow6 = (~(Y67ow6 & F77ow6));
assign F77ow6 = (M77ow6 & T77ow6);
assign T77ow6 = (A87ow6 & H87ow6);
assign H87ow6 = (~(O87ow6 & V87ow6));
assign V87ow6 = (~(Q1ziu6 | Gaziu6));
assign Q1ziu6 = (!Y31ju6);
assign O87ow6 = (Nyiiu6 & Evyiu6);
assign A87ow6 = (~(Ipziu6 & S6aiu6));
assign Ipziu6 = (~(Lkaiu6 | Dxziu6));
assign M77ow6 = (C97ow6 & J97ow6);
assign J97ow6 = (~(Q97ow6 & X97ow6));
assign C97ow6 = (~(Vviiu6 & Ea7ow6));
assign Ea7ow6 = (~(Nj6ow6 & La7ow6));
assign La7ow6 = (~(Y40ju6 & Db0ju6));
assign Y67ow6 = (Sa7ow6 & Za7ow6);
assign Za7ow6 = (Kgaiu6 | Wthiu6);
assign Wthiu6 = (!K2aiu6);
assign Sa7ow6 = (Gb7ow6 & Nb7ow6);
assign Nb7ow6 = (~(Ub7ow6 & Q5aiu6));
assign Ub7ow6 = (~(Bc7ow6 & Ic7ow6));
assign Ic7ow6 = (~(Pc7ow6 & Wc7ow6));
assign Wc7ow6 = (~(H95iu6 | Oviiu6));
assign Pc7ow6 = (Dmiiu6 & Jwiiu6);
assign Bc7ow6 = (~(Dd7ow6 & J8ziu6));
assign J8ziu6 = (Kd7ow6 & Wh0ju6);
assign Kd7ow6 = (~(Ph0ju6 | D7fpw6[5]));
assign Ph0ju6 = (Aq1ju6 | D7fpw6[7]);
assign Gb7ow6 = (~(Uyiiu6 & Rd7ow6));
assign Rd7ow6 = (~(Yd7ow6 & Fe7ow6));
assign Fe7ow6 = (~(Wliiu6 & Me7ow6));
assign Me7ow6 = (~(Ftjiu6 & Te7ow6));
assign Te7ow6 = (~(Af7ow6 & Uriiu6));
assign Af7ow6 = (~(Hf7ow6 & Of7ow6));
assign Of7ow6 = (Vf7ow6 & Cg7ow6);
assign Cg7ow6 = (Ar0ju6 | D7fpw6[10]);
assign Vf7ow6 = (Hk0ju6 | Kcziu6);
assign Hf7ow6 = (Qz0ju6 & D7fpw6[14]);
assign Qz0ju6 = (Jg7ow6 & Qg7ow6);
assign Qg7ow6 = (~(Xg7ow6 & D7fpw6[7]));
assign Jg7ow6 = (~(D7fpw6[10] & Eh7ow6));
assign Eh7ow6 = (D7fpw6[8] | Qe0ju6);
assign Qe0ju6 = (!Rg2ju6);
assign Yd7ow6 = (~(Dmiiu6 & Lh7ow6));
assign Lh7ow6 = (~(Sh7ow6 & Zh7ow6));
assign Zh7ow6 = (H95iu6 | D7fpw6[9]);
assign Sh7ow6 = (Z01ju6 & Gi7ow6);
assign Gi7ow6 = (Wiliu6 | Gaziu6);
assign Z01ju6 = (~(Qxoiu6 & Nbkiu6));
assign J27ow6 = (Ni7ow6 & K0jiu6);
assign Ni7ow6 = (Ui7ow6 & Bj7ow6);
assign Bj7ow6 = (~(Moaiu6 & Us2ju6));
assign Ui7ow6 = (Qojiu6 | Cyfpw6[7]);
assign Ssohu6 = (Ij7ow6 | Pj7ow6);
assign Pj7ow6 = (~(Wj7ow6 | Dk7ow6));
assign Ij7ow6 = (Rk7ow6 ? S8fpw6[5] : Kk7ow6);
assign Kk7ow6 = (~(Yk7ow6 & Fl7ow6));
assign Fl7ow6 = (Ml7ow6 & Tl7ow6);
assign Tl7ow6 = (~(Am7ow6 & Ppfpw6[5]));
assign Ml7ow6 = (Dzjiu6 | Hm7ow6);
assign Yk7ow6 = (Om7ow6 & Vm7ow6);
assign Vm7ow6 = (~(Cbbiu6 & D7fpw6[10]));
assign Om7ow6 = (A1kiu6 | Cn7ow6);
assign Lsohu6 = (O25iu6 ? X3fpw6[0] : Jn7ow6);
assign O25iu6 = (~(HREADY & Qn7ow6));
assign Qn7ow6 = (~(Xn7ow6 & Eo7ow6));
assign Eo7ow6 = (Lo7ow6 & So7ow6);
assign So7ow6 = (~(Zo7ow6 | Ujjiu6));
assign Zo7ow6 = (~(Isiiu6 & Dz6ow6));
assign Isiiu6 = (~(Gp7ow6 & Np7ow6));
assign Np7ow6 = (~(Xe8iu6 | Cyfpw6[4]));
assign Gp7ow6 = (~(R2aiu6 | Xojiu6));
assign Lo7ow6 = (Up7ow6 & Bq7ow6);
assign Bq7ow6 = (~(Iq7ow6 & Cyfpw6[0]));
assign Iq7ow6 = (~(Kq0iu6 | Cyfpw6[3]));
assign Up7ow6 = (Pq7ow6 & Wq7ow6);
assign Wq7ow6 = (~(Dr7ow6 & Kr7ow6));
assign Dr7ow6 = (L45iu6 & Zraiu6);
assign Pq7ow6 = (~(Rr7ow6 & Y31ju6));
assign Rr7ow6 = (M7kiu6 & Yr7ow6);
assign Yr7ow6 = (D7fpw6[14] | Fs7ow6);
assign Xn7ow6 = (Ms7ow6 & Ts7ow6);
assign Ts7ow6 = (At7ow6 & Ht7ow6);
assign Ht7ow6 = (~(Ot7ow6 & D7fpw6[3]));
assign At7ow6 = (Vt7ow6 & Cu7ow6);
assign Cu7ow6 = (~(Zzniu6 & Ju7ow6));
assign Ju7ow6 = (Qu7ow6 | Ae0iu6);
assign Vt7ow6 = (~(U98iu6 & Xu7ow6));
assign Xu7ow6 = (Mo2ju6 | Us2ju6);
assign Ms7ow6 = (Ev7ow6 & Lv7ow6);
assign Ev7ow6 = (Sv7ow6 & Zv7ow6);
assign Zv7ow6 = (~(Uyiiu6 & Gw7ow6));
assign Gw7ow6 = (~(Nw7ow6 & Uw7ow6));
assign Uw7ow6 = (~(Bx7ow6 & Dmiiu6));
assign Bx7ow6 = (Nbkiu6 & Zraiu6);
assign Nw7ow6 = (Ix7ow6 & Px7ow6);
assign Px7ow6 = (~(Wx7ow6 & Dy7ow6));
assign Dy7ow6 = (Ky7ow6 & Ry7ow6);
assign Ky7ow6 = (L88iu6 & Dzjiu6);
assign L88iu6 = (~(Ndiiu6 | Gkiiu6));
assign Wx7ow6 = (~(Kcziu6 | U5jiu6));
assign Ix7ow6 = (~(Yy7ow6 & Fz7ow6));
assign Fz7ow6 = (Th2ju6 & Ak0ju6);
assign Yy7ow6 = (Cwiiu6 & Aujiu6);
assign Sv7ow6 = (~(Y0jiu6 & Gwyiu6));
assign Jn7ow6 = (~(Mz7ow6 & Tz7ow6));
assign Tz7ow6 = (A08ow6 & H08ow6);
assign H08ow6 = (R75iu6 | I65iu6);
assign I65iu6 = (!S8fpw6[8]);
assign A08ow6 = (O08ow6 & V08ow6);
assign V08ow6 = (~(L45iu6 & C18ow6));
assign C18ow6 = (~(J18ow6 & Q18ow6));
assign Q18ow6 = (X18ow6 & E28ow6);
assign E28ow6 = (L28ow6 | Eoyiu6);
assign X18ow6 = (~(Zoyiu6 & G55iu6));
assign J18ow6 = (S28ow6 & Z28ow6);
assign Z28ow6 = (B65iu6 | N55iu6);
assign S28ow6 = (P65iu6 | S8fpw6[8]);
assign P65iu6 = (!S8fpw6[9]);
assign O08ow6 = (~(D7fpw6[3] & K75iu6));
assign K75iu6 = (~(Wiliu6 & G38ow6));
assign G38ow6 = (N38ow6 | I6jiu6);
assign Mz7ow6 = (U38ow6 & Gpyiu6);
assign Gpyiu6 = (B48ow6 & F85iu6);
assign F85iu6 = (K0jiu6 & Twniu6);
assign K0jiu6 = (R2aiu6 | Tr0iu6);
assign B48ow6 = (~(N20ju6 | Hzziu6));
assign U38ow6 = (I48ow6 & P48ow6);
assign P48ow6 = (~(A95iu6 & D7fpw6[0]));
assign I48ow6 = (H95iu6 | Ad8iu6);
assign Esohu6 = (~(W48ow6 & D58ow6));
assign D58ow6 = (K58ow6 & R58ow6);
assign R58ow6 = (~(Egziu6 & Eafpw6[7]));
assign K58ow6 = (Y58ow6 & Sgziu6);
assign Y58ow6 = (~(Zgziu6 & Qukiu6));
assign Qukiu6 = (~(F68ow6 & M68ow6));
assign M68ow6 = (T68ow6 & A78ow6);
assign A78ow6 = (Cfliu6 | H78ow6);
assign T68ow6 = (O78ow6 & Mdliu6);
assign O78ow6 = (~(Qfliu6 & V78ow6));
assign F68ow6 = (C88ow6 & J88ow6);
assign J88ow6 = (Ycliu6 | Q88ow6);
assign C88ow6 = (~(Aeliu6 & X88ow6));
assign W48ow6 = (E98ow6 & L98ow6);
assign L98ow6 = (~(Zsfpw6[6] & Cmziu6));
assign E98ow6 = (~(vis_pc_o[6] & Jmziu6));
assign Xrohu6 = (~(S98ow6 & Z98ow6));
assign Z98ow6 = (Ga8ow6 & Na8ow6);
assign Na8ow6 = (~(Egziu6 & Eafpw6[31]));
assign Ga8ow6 = (Ua8ow6 & Sgziu6);
assign Ua8ow6 = (Ft6ow6 | Ualiu6);
assign Ualiu6 = (Bb8ow6 & Ib8ow6);
assign Ib8ow6 = (Pb8ow6 & Wb8ow6);
assign Wb8ow6 = (~(Dc8ow6 & X88ow6));
assign Pb8ow6 = (Kc8ow6 & Djziu6);
assign Kc8ow6 = (~(Rc8ow6 & V78ow6));
assign Bb8ow6 = (Yc8ow6 & Fd8ow6);
assign Fd8ow6 = (Mkziu6 | Q88ow6);
assign Yc8ow6 = (Hlziu6 | H78ow6);
assign S98ow6 = (Md8ow6 & Td8ow6);
assign Td8ow6 = (~(Zsfpw6[30] & Cmziu6));
assign Md8ow6 = (~(vis_pc_o[30] & Jmziu6));
assign Qrohu6 = (Ae8ow6 | He8ow6);
assign He8ow6 = (~(Oe8ow6 | Cyfpw6[6]));
assign Ae8ow6 = (HREADY ? Ve8ow6 : Cyfpw6[1]);
assign Ve8ow6 = (~(Cf8ow6 & Jf8ow6));
assign Jf8ow6 = (Qf8ow6 & Xf8ow6);
assign Xf8ow6 = (Eg8ow6 & Lg8ow6);
assign Lg8ow6 = (~(Sg8ow6 & Neoiu6));
assign Sg8ow6 = (Zg8ow6 & Mr0iu6);
assign Zg8ow6 = (~(E4jiu6 & Gh8ow6));
assign Gh8ow6 = (~(Nh8ow6 & Pthiu6));
assign Nh8ow6 = (~(R75iu6 | Cyfpw6[5]));
assign Eg8ow6 = (~(Uh8ow6 & Hiaiu6));
assign Uh8ow6 = (Bi8ow6 & Q5aiu6);
assign Bi8ow6 = (~(Ii8ow6 & Pi8ow6));
assign Pi8ow6 = (Wi8ow6 & Dj8ow6);
assign Dj8ow6 = (~(J9kiu6 & Kj8ow6));
assign Kj8ow6 = (~(Rj8ow6 & Yj8ow6));
assign Yj8ow6 = (Fk8ow6 & S01ju6);
assign S01ju6 = (!Fs7ow6);
assign Fs7ow6 = (D7fpw6[11] & I6jiu6);
assign Fk8ow6 = (~(Mk8ow6 & X1ziu6));
assign Mk8ow6 = (Zwciu6 | D7fpw6[8]);
assign Zwciu6 = (!Jehhu6);
assign Rj8ow6 = (Tk8ow6 & Al8ow6);
assign Al8ow6 = (Hl8ow6 | D7fpw6[11]);
assign Tk8ow6 = (D7fpw6[13] | D7fpw6[8]);
assign Wi8ow6 = (Ol8ow6 & Vl8ow6);
assign Vl8ow6 = (~(Cm8ow6 & Jm8ow6));
assign Jm8ow6 = (~(I6jiu6 | Jjhiu6));
assign Cm8ow6 = (Y40ju6 & Nyiiu6);
assign Nyiiu6 = (D7fpw6[11] & Ftjiu6);
assign Ol8ow6 = (~(Qm8ow6 & Evyiu6));
assign Qm8ow6 = (~(Oviiu6 | Gaziu6));
assign Ii8ow6 = (~(Xm8ow6 | En8ow6));
assign En8ow6 = (Ejiiu6 & Dmiiu6);
assign Dmiiu6 = (Jiiiu6 & D7fpw6[14]);
assign Xm8ow6 = (S1ehu6 ? Sn8ow6 : Ln8ow6);
assign Ln8ow6 = (~(Zn8ow6 & Go8ow6));
assign Go8ow6 = (No8ow6 | Lroiu6);
assign Lroiu6 = (!Ejiiu6);
assign No8ow6 = (!Il3ju6);
assign Zn8ow6 = (Uo8ow6 & Xs0ju6);
assign Xs0ju6 = (Wiliu6 | Co6ow6);
assign Wiliu6 = (!Mtjiu6);
assign Uo8ow6 = (~(Bp8ow6 & Mtjiu6));
assign Bp8ow6 = (D7fpw6[14] & Ip8ow6);
assign Ip8ow6 = (~(Pp8ow6 & Wp8ow6));
assign Wp8ow6 = (Aq1ju6 ? Dq8ow6 : D7fpw6[9]);
assign Aq1ju6 = (~(D7fpw6[8] & Ad8iu6));
assign Dq8ow6 = (U5jiu6 | O95iu6);
assign Pp8ow6 = (Kq8ow6 & Oviiu6);
assign Kq8ow6 = (~(D7fpw6[8] & Rq8ow6));
assign Rq8ow6 = (~(Yq8ow6 & Fr8ow6));
assign Fr8ow6 = (I6jiu6 | D7fpw6[7]);
assign Yq8ow6 = (~(Db0ju6 | Dcziu6));
assign Qf8ow6 = (Mr8ow6 & Tr8ow6);
assign Tr8ow6 = (~(As8ow6 & Hs8ow6));
assign As8ow6 = (Frziu6 & Hzziu6);
assign Mr8ow6 = (~(Os8ow6 & Geaiu6));
assign Os8ow6 = (~(Vs8ow6 & Ct8ow6));
assign Ct8ow6 = (~(Jt8ow6 & Vs0iu6));
assign Vs0iu6 = (F86ow6 & Cyfpw6[0]);
assign F86ow6 = (~(Knaiu6 | Tfjiu6));
assign Jt8ow6 = (Qe8iu6 & Gwyiu6);
assign Vs8ow6 = (~(Qt8ow6 & D7fpw6[11]));
assign Qt8ow6 = (Xt8ow6 & Q5aiu6);
assign Xt8ow6 = (Ry7ow6 | Zakiu6);
assign Zakiu6 = (Th2ju6 & I6jiu6);
assign Ry7ow6 = (!Oaiiu6);
assign Cf8ow6 = (Eu8ow6 & Lu8ow6);
assign Lu8ow6 = (Su8ow6 & Zu8ow6);
assign Zu8ow6 = (~(Gv8ow6 & Zraiu6));
assign Gv8ow6 = (~(Nv8ow6 & Uv8ow6));
assign Uv8ow6 = (Bw8ow6 & Td0iu6);
assign Bw8ow6 = (Re6ow6 & Iw8ow6);
assign Re6ow6 = (~(Pw8ow6 & Ww8ow6));
assign Pw8ow6 = (~(Iuniu6 | Xmliu6));
assign Nv8ow6 = (Dx8ow6 & Kx8ow6);
assign Kx8ow6 = (~(U0aiu6 & Rx8ow6));
assign Rx8ow6 = (Tfjiu6 | X97ow6);
assign Dx8ow6 = (~(S6aiu6 & Yx8ow6));
assign Yx8ow6 = (Geoiu6 | Ly2ju6);
assign Ly2ju6 = (Vo3ju6 & Tr0iu6);
assign Eu8ow6 = (Fy8ow6 & My8ow6);
assign My8ow6 = (Ty8ow6 | Xe8iu6);
assign Fy8ow6 = (Dxziu6 ? Hz8ow6 : Az8ow6);
assign Hz8ow6 = (~(Oz8ow6 & Moaiu6));
assign Oz8ow6 = (Toaiu6 & Cyfpw6[7]);
assign Az8ow6 = (~(Vz8ow6 & F9aju6));
assign Vz8ow6 = (Ls1ju6 & Sq3ju6);
assign Jrohu6 = (C09ow6 & J09ow6);
assign J09ow6 = (~(Q09ow6 & X09ow6));
assign X09ow6 = (E19ow6 & L19ow6);
assign L19ow6 = (S19ow6 & Z19ow6);
assign Z19ow6 = (G29ow6 & Yryiu6);
assign Yryiu6 = (~(Ujjiu6 & Bkjiu6));
assign G29ow6 = (~(N29ow6 & Cyfpw6[0]));
assign N29ow6 = (U29ow6 & B39ow6);
assign B39ow6 = (~(I39ow6 & R75iu6));
assign I39ow6 = (~(P39ow6 & Yljiu6));
assign P39ow6 = (~(Hs0iu6 | Dxziu6));
assign U29ow6 = (Difiu6 | Pugiu6);
assign Difiu6 = (Cyfpw6[6] & Ii0iu6);
assign S19ow6 = (W39ow6 & D49ow6);
assign D49ow6 = (~(K49ow6 & T23ju6));
assign K49ow6 = (~(C0ehu6 | Cyfpw6[7]));
assign W39ow6 = (~(R49ow6 & W0piu6));
assign R49ow6 = (D7fpw6[11] & Y49ow6);
assign Y49ow6 = (~(C27ow6 & F59ow6));
assign F59ow6 = (~(M59ow6 & C0ehu6));
assign M59ow6 = (~(X1ziu6 | D7fpw6[10]));
assign E19ow6 = (T59ow6 & A69ow6);
assign A69ow6 = (H69ow6 & O69ow6);
assign O69ow6 = (~(V69ow6 & Hzziu6));
assign V69ow6 = (~(Yp8iu6 | Y7ghu6));
assign H69ow6 = (~(C79ow6 & J79ow6));
assign C79ow6 = (Yljiu6 & Taaiu6);
assign T59ow6 = (Q79ow6 & X79ow6);
assign X79ow6 = (~(Hwaiu6 & A3aju6));
assign Hwaiu6 = (~(R75iu6 | Knaiu6));
assign Q79ow6 = (~(Dxziu6 & E89ow6));
assign E89ow6 = (~(L89ow6 & S89ow6));
assign S89ow6 = (~(Z89ow6 & X97ow6));
assign Z89ow6 = (D1piu6 & Tfjiu6);
assign L89ow6 = (~(Jf6ju6 & N3ziu6));
assign Q09ow6 = (G99ow6 & N99ow6);
assign N99ow6 = (U99ow6 & Ba9ow6);
assign Ba9ow6 = (Ia9ow6 & Pa9ow6);
assign Pa9ow6 = (~(Uyiiu6 & Wa9ow6));
assign Wa9ow6 = (~(Xl0ju6 & Db9ow6));
assign Db9ow6 = (~(Kb9ow6 & Ftjiu6));
assign Kb9ow6 = (~(Biliu6 & Rb9ow6));
assign Rb9ow6 = (Yb9ow6 | I6jiu6);
assign Biliu6 = (!Sn8ow6);
assign Sn8ow6 = (C0ehu6 & X1ziu6);
assign Ia9ow6 = (Thaiu6 | Cyfpw6[5]);
assign U99ow6 = (Fc9ow6 & Mc9ow6);
assign Mc9ow6 = (~(De6ow6 & Vxniu6));
assign Fc9ow6 = (Iw8ow6 | Ae0iu6);
assign G99ow6 = (Tc9ow6 & Ad9ow6);
assign Ad9ow6 = (Hd9ow6 & Od9ow6);
assign Od9ow6 = (~(S6aiu6 & Vd9ow6));
assign Vd9ow6 = (~(Ce9ow6 & Je9ow6));
assign Je9ow6 = (Nlaiu6 ? Ey2ju6 : Cyfpw6[1]);
assign Ce9ow6 = (~(Qe9ow6 | Ep6ow6));
assign Qe9ow6 = (~(Lkaiu6 | Eoyiu6));
assign Hd9ow6 = (Xe9ow6 | Wxyiu6);
assign Wxyiu6 = (L62ju6 & Zraiu6);
assign L62ju6 = (!Nsaiu6);
assign Tc9ow6 = (T41ju6 & Ef9ow6);
assign Ef9ow6 = (~(Lf9ow6 & Q5aiu6));
assign Lf9ow6 = (~(Sf9ow6 & Zf9ow6));
assign Zf9ow6 = (Gg9ow6 & Ng9ow6);
assign Ng9ow6 = (~(Ug9ow6 & Vboiu6));
assign Ug9ow6 = (~(R75iu6 | H4ghu6));
assign Gg9ow6 = (Bh9ow6 & Ih9ow6);
assign Ih9ow6 = (~(Ph9ow6 & P0piu6));
assign Ph9ow6 = (Wh9ow6 & Ftjiu6);
assign Wh9ow6 = (Di9ow6 | Ki9ow6);
assign Ki9ow6 = (Tniiu6 ? Dcziu6 : Ad8iu6);
assign Di9ow6 = (~(Ri9ow6 & Ar0ju6));
assign Ar0ju6 = (!Jz0ju6);
assign Ri9ow6 = (Ndiiu6 | O95iu6);
assign Bh9ow6 = (~(Yi9ow6 & Db0ju6));
assign Yi9ow6 = (~(H95iu6 | X1ziu6));
assign H95iu6 = (!Ozziu6);
assign Sf9ow6 = (Fj9ow6 & Mj9ow6);
assign Mj9ow6 = (~(Xiiiu6 & Tj9ow6));
assign Tj9ow6 = (~(Ak9ow6 & Hk9ow6));
assign Hk9ow6 = (~(Aujiu6 & U5jiu6));
assign U5jiu6 = (!Jwiiu6);
assign Ak9ow6 = (~(Ok9ow6 | Vk9ow6));
assign Ok9ow6 = (Y40ju6 & Cl9ow6);
assign Cl9ow6 = (~(Jl9ow6 & Ql9ow6));
assign Ql9ow6 = (Oviiu6 | D7fpw6[6]);
assign Jl9ow6 = (~(Dcziu6 | D7fpw6[8]));
assign Fj9ow6 = (Xl9ow6 & Em9ow6);
assign Em9ow6 = (~(Hl8ow6 & Lm9ow6));
assign Lm9ow6 = (~(S80ju6 & Sm9ow6));
assign Sm9ow6 = (~(J9kiu6 & Zm9ow6));
assign Zm9ow6 = (~(Gn9ow6 & Nn9ow6));
assign Nn9ow6 = (Un9ow6 & I6jiu6);
assign Un9ow6 = (D7fpw6[4] | D7fpw6[6]);
assign Gn9ow6 = (~(O95iu6 | Dzjiu6));
assign Xl9ow6 = (~(C0ehu6 & Bo9ow6));
assign Bo9ow6 = (~(Io9ow6 & Po9ow6));
assign Po9ow6 = (~(Wo9ow6 & Aujiu6));
assign Wo9ow6 = (~(X1ziu6 | D7fpw6[8]));
assign Io9ow6 = (Dp9ow6 & Uriiu6);
assign Dp9ow6 = (~(Kp9ow6 & Y40ju6));
assign Kp9ow6 = (~(Jwiiu6 | D7fpw6[15]));
assign T41ju6 = (Rp9ow6 & Yp9ow6);
assign Yp9ow6 = (Fq9ow6 & B1aiu6);
assign Fq9ow6 = (~(Mq9ow6 & Cyfpw6[4]));
assign Mq9ow6 = (~(Geaiu6 | Cyfpw6[5]));
assign Rp9ow6 = (HREADY & Tq9ow6);
assign C09ow6 = (Cyfpw6[0] | HREADY);
assign Crohu6 = (Ar9ow6 & Hr9ow6);
assign Hr9ow6 = (~(Or9ow6 & Vr9ow6));
assign Vr9ow6 = (Cs9ow6 & Js9ow6);
assign Js9ow6 = (Qs9ow6 & Xs9ow6);
assign Xs9ow6 = (Et9ow6 & A42ju6);
assign A42ju6 = (~(Lt9ow6 & Htyiu6));
assign Lt9ow6 = (Th2ju6 & St9ow6);
assign St9ow6 = (~(D7fpw6[12] & Zt9ow6));
assign Et9ow6 = (~(Ujjiu6 | Ot7ow6));
assign Ot7ow6 = (Gu9ow6 & Nu9ow6);
assign Gu9ow6 = (~(Jcaiu6 | Cyfpw6[0]));
assign Ujjiu6 = (Uu9ow6 & D7fpw6[15]);
assign Qs9ow6 = (Bv9ow6 & Iv9ow6);
assign Iv9ow6 = (~(Pv9ow6 & Wv9ow6));
assign Wv9ow6 = (D7fpw6[11] & Dw9ow6);
assign Dw9ow6 = (Gkiiu6 | Fp1ju6);
assign Pv9ow6 = (Yv1ju6 & Nbkiu6);
assign Bv9ow6 = (~(Kw9ow6 & Rw9ow6));
assign Rw9ow6 = (~(D7fpw6[5] | D7fpw6[7]));
assign Kw9ow6 = (~(P82ju6 | Yw9ow6));
assign Yw9ow6 = (D7fpw6[4] & D7fpw6[6]);
assign Cs9ow6 = (Fx9ow6 & Mx9ow6);
assign Mx9ow6 = (Tx9ow6 & Ay9ow6);
assign Ay9ow6 = (~(Hy9ow6 & Vviiu6));
assign Hy9ow6 = (Hiaiu6 & Oy9ow6);
assign Oy9ow6 = (~(Vy9ow6 & Cz9ow6));
assign Cz9ow6 = (Jz9ow6 | Gaziu6);
assign Vy9ow6 = (X1ziu6 | Gkiiu6);
assign Tx9ow6 = (~(Qz9ow6 & Htyiu6));
assign Qz9ow6 = (Xz9ow6 & Zraiu6);
assign Xz9ow6 = (~(E0aow6 & L0aow6));
assign L0aow6 = (~(X8ziu6 & A95iu6));
assign X8ziu6 = (~(D7fpw6[11] | D7fpw6[8]));
assign E0aow6 = (S80ju6 | Gaziu6);
assign Fx9ow6 = (S0aow6 & Z0aow6);
assign Z0aow6 = (~(G1aow6 & K2aiu6));
assign G1aow6 = (N1aow6 & Y2oiu6);
assign S0aow6 = (~(U1aow6 & Neoiu6));
assign U1aow6 = (Omyiu6 & B2aow6);
assign B2aow6 = (~(I2aow6 & P2aow6));
assign P2aow6 = (Vwaiu6 | Mr0iu6);
assign I2aow6 = (~(G47ow6 | W2aow6));
assign Or9ow6 = (D3aow6 & K3aow6);
assign K3aow6 = (R3aow6 & Y3aow6);
assign Y3aow6 = (F4aow6 & M4aow6);
assign M4aow6 = (Tdziu6 | Qpaju6);
assign Tdziu6 = (~(Q97ow6 & T4aow6));
assign Q97ow6 = (~(E4jiu6 | Cyfpw6[0]));
assign F4aow6 = (A5aow6 & H5aow6);
assign H5aow6 = (~(O5aow6 & Yo1ju6));
assign O5aow6 = (D7fpw6[14] & V5aow6);
assign V5aow6 = (C6aow6 | J6aow6);
assign J6aow6 = (D7fpw6[7] ? X6aow6 : Q6aow6);
assign X6aow6 = (~(Jz0ju6 | D7fpw6[10]));
assign Jz0ju6 = (Ad8iu6 & Ndiiu6);
assign C6aow6 = (~(E7aow6 & Hk0ju6));
assign Hk0ju6 = (!Fp1ju6);
assign Fp1ju6 = (I6jiu6 & Tniiu6);
assign E7aow6 = (L7aow6 | D7fpw6[9]);
assign A5aow6 = (~(Pthiu6 & S7aow6));
assign S7aow6 = (~(Z7aow6 & G8aow6));
assign G8aow6 = (Jojiu6 | Y2oiu6);
assign Z7aow6 = (~(Ls1ju6 & Cyfpw6[5]));
assign R3aow6 = (N8aow6 & U8aow6);
assign U8aow6 = (~(B9aow6 & Geaiu6));
assign B9aow6 = (~(I9aow6 & P9aow6));
assign P9aow6 = (R2aiu6 | Y2oiu6);
assign I9aow6 = (W9aow6 & Daaow6);
assign Daaow6 = (~(Kaaow6 & Raaow6));
assign Kaaow6 = (M7kiu6 & X1ziu6);
assign M7kiu6 = (Yaaow6 & Ozziu6);
assign Yaaow6 = (~(Ae0iu6 | D7fpw6[15]));
assign W9aow6 = (Jxoiu6 | Ak0ju6);
assign Ak0ju6 = (Qxoiu6 & Ndiiu6);
assign Jxoiu6 = (~(Fbaow6 & R7jiu6));
assign Fbaow6 = (Ia8iu6 & Q5aiu6);
assign N8aow6 = (~(Dxziu6 & Mbaow6));
assign Mbaow6 = (~(Tbaow6 & Acaow6));
assign Acaow6 = (~(Ls1ju6 & Hcaow6));
assign Hcaow6 = (Rljiu6 | Ocaow6);
assign Ocaow6 = (~(Qjaiu6 | Cyfpw6[0]));
assign Tbaow6 = (Vcaow6 & Cdaow6);
assign Cdaow6 = (~(Jdaow6 & Qdaow6));
assign Qdaow6 = (Qe8iu6 & Mr0iu6);
assign Jdaow6 = (Eoyiu6 & Geoiu6);
assign Geoiu6 = (Wp0iu6 & Ii0iu6);
assign Eoyiu6 = (~(L28ow6 | S8fpw6[7]));
assign Vcaow6 = (~(Xdaow6 & Vxniu6));
assign Xdaow6 = (D1piu6 & Zraiu6);
assign D3aow6 = (Eeaow6 & Leaow6);
assign Leaow6 = (Seaow6 & Zeaow6);
assign Zeaow6 = (~(Hs8ow6 & Nriiu6));
assign Seaow6 = (Qojiu6 | M32ju6);
assign Qojiu6 = (!M2piu6);
assign Eeaow6 = (Ez1ju6 & Oeziu6);
assign Oeziu6 = (Gfaow6 & HREADY);
assign Gfaow6 = (Thaiu6 & Dz6ow6);
assign Thaiu6 = (E45iu6 | Y2oiu6);
assign Ez1ju6 = (Nfaow6 & J5aiu6);
assign J5aiu6 = (Qp3ju6 | Jojiu6);
assign Qp3ju6 = (!J79ow6);
assign Nfaow6 = (Ufaow6 & Bgaow6);
assign Ufaow6 = (H3piu6 | Cyfpw6[6]);
assign H3piu6 = (!C78iu6);
assign C78iu6 = (S6aiu6 & Neoiu6);
assign Ar9ow6 = (Cyfpw6[4] | HREADY);
assign Vqohu6 = (!Igaow6);
assign Igaow6 = (HREADY ? Pgaow6 : Xe8iu6);
assign Pgaow6 = (Wgaow6 & Dhaow6);
assign Dhaow6 = (Khaow6 & Rhaow6);
assign Rhaow6 = (Yhaow6 & Fiaow6);
assign Fiaow6 = (Miaow6 & Tiaow6);
assign Tiaow6 = (~(Ajaow6 & Hjaow6));
assign Hjaow6 = (~(Qpaju6 | D7fpw6[13]));
assign Ajaow6 = (Raaow6 & Imaiu6);
assign Miaow6 = (Imoiu6 & Dz6ow6);
assign Dz6ow6 = (~(Ojaow6 & N20ju6));
assign Ojaow6 = (~(Ii0iu6 | Lraiu6));
assign Imoiu6 = (~(Pfoiu6 & Pu1ju6));
assign Yhaow6 = (Vjaow6 & Ckaow6);
assign Ckaow6 = (~(Jkaow6 & Qkaow6));
assign Qkaow6 = (L45iu6 & Oiaiu6);
assign Jkaow6 = (~(Wfoiu6 | Xkaow6));
assign Vjaow6 = (~(Elaow6 & J79ow6));
assign Elaow6 = (U98iu6 & Taaiu6);
assign U98iu6 = (Llaow6 & Jjhiu6);
assign Khaow6 = (Slaow6 & Zlaow6);
assign Zlaow6 = (Gmaow6 & Nmaow6);
assign Nmaow6 = (~(Llaow6 & Umaow6));
assign Umaow6 = (~(Bnaow6 & Inaow6));
assign Inaow6 = (~(Pnaow6 & Ruaiu6));
assign Pnaow6 = (~(Wnaow6 & Doaow6));
assign Doaow6 = (Koaow6 & Xa6ow6);
assign Xa6ow6 = (~(Roaow6 & Cyfpw6[7]));
assign Roaow6 = (~(Geaiu6 | Cyfpw6[3]));
assign Koaow6 = (~(Yoaow6 & Hzziu6));
assign Yoaow6 = (Fpaow6 & Mr0iu6);
assign Fpaow6 = (~(Mpaow6 & Tpaow6));
assign Tpaow6 = (X1ziu6 | S1ehu6);
assign Wnaow6 = (Aqaow6 & Hqaow6);
assign Hqaow6 = (Z6oiu6 | Geaiu6);
assign Aqaow6 = (R75iu6 | Cyfpw6[6]);
assign Bnaow6 = (~(Nu9ow6 & V4aiu6));
assign Gmaow6 = (Oqaow6 & Vqaow6);
assign Vqaow6 = (~(Yi7ju6 & Pu1ju6));
assign Yi7ju6 = (~(Ii0iu6 | Cyfpw6[6]));
assign Oqaow6 = (~(Yo1ju6 & Craow6));
assign Craow6 = (~(Jraow6 & Qraow6));
assign Qraow6 = (L7aow6 | O7ziu6);
assign Jraow6 = (~(D7fpw6[8] & Xraow6));
assign Xraow6 = (~(Esaow6 & Lsaow6));
assign Lsaow6 = (~(D7fpw6[9] & Dcziu6));
assign Esaow6 = (~(Qxoiu6 & O95iu6));
assign Yo1ju6 = (Ba8iu6 & Ssaow6);
assign Ba8iu6 = (~(S80ju6 | D7fpw6[13]));
assign Slaow6 = (Zsaow6 & Gtaow6);
assign Gtaow6 = (~(Ntaow6 & Zraiu6));
assign Ntaow6 = (~(Rz6ow6 & Utaow6));
assign Utaow6 = (Gtgiu6 | Iuniu6);
assign Gtgiu6 = (!Buaow6);
assign Rz6ow6 = (~(Iuaow6 & Nu9ow6));
assign Iuaow6 = (~(Nlaiu6 | H4ghu6));
assign Zsaow6 = (~(Rljiu6 & It2ju6));
assign Rljiu6 = (Xzmiu6 & Cyfpw6[5]);
assign Wgaow6 = (Puaow6 & Wuaow6);
assign Wuaow6 = (Dvaow6 & Kvaow6);
assign Kvaow6 = (Rvaow6 & Yvaow6);
assign Yvaow6 = (Rb0ju6 | Fwaow6);
assign Rb0ju6 = (~(Bziiu6 & Oviiu6));
assign Rvaow6 = (Mwaow6 & Twaow6);
assign Twaow6 = (~(D7fpw6[12] & Axaow6));
assign Axaow6 = (~(Hxaow6 & Oxaow6));
assign Oxaow6 = (Fwaow6 | N38ow6);
assign Fwaow6 = (!Ssaow6);
assign Hxaow6 = (Vxaow6 & Cyaow6);
assign Cyaow6 = (~(Jyaow6 & Qyaow6));
assign Qyaow6 = (Xyaow6 & Geaiu6);
assign Xyaow6 = (~(Jz9ow6 & Ezaow6));
assign Ezaow6 = (O7ziu6 | Ndiiu6);
assign Jz9ow6 = (~(Xg7ow6 & Cwiiu6));
assign Xg7ow6 = (~(Tniiu6 | D7fpw6[8]));
assign Jyaow6 = (Vviiu6 & Kxziu6);
assign Vxaow6 = (~(Lzaow6 & W82ju6));
assign W82ju6 = (Szaow6 & D7fpw6[5]);
assign Szaow6 = (~(D7fpw6[6] | D7fpw6[7]));
assign Lzaow6 = (~(P82ju6 | A1kiu6));
assign P82ju6 = (~(Zzaow6 & G0bow6));
assign G0bow6 = (Rmiiu6 & D7fpw6[8]);
assign Rmiiu6 = (F6ziu6 & Th2ju6);
assign Zzaow6 = (Wh0ju6 & Htyiu6);
assign Mwaow6 = (~(Hzziu6 & N0bow6));
assign N0bow6 = (~(U0bow6 & B1bow6));
assign B1bow6 = (~(Oxniu6 & Tfjiu6));
assign U0bow6 = (I1bow6 & P1bow6);
assign I1bow6 = (~(W1bow6 & Ia8iu6));
assign W1bow6 = (Aujiu6 & Frziu6);
assign Dvaow6 = (D2bow6 & K2bow6);
assign K2bow6 = (~(Qe8iu6 & R2bow6));
assign R2bow6 = (~(Y2bow6 & F3bow6));
assign F3bow6 = (~(J79ow6 | D31ju6));
assign Y2bow6 = (M3bow6 & T3bow6);
assign T3bow6 = (Jc2ju6 | Knaiu6);
assign M3bow6 = (~(Frziu6 & K2aiu6));
assign D2bow6 = (~(D7fpw6[11] & A4bow6));
assign A4bow6 = (~(H4bow6 & O4bow6));
assign O4bow6 = (V4bow6 & C5bow6);
assign C5bow6 = (~(J5bow6 & Yv1ju6));
assign Yv1ju6 = (Ssaow6 & X1ziu6);
assign J5bow6 = (~(Tniiu6 | Jjhiu6));
assign V4bow6 = (~(Q5bow6 & Htyiu6));
assign Q5bow6 = (~(C27ow6 | Ae0iu6));
assign H4bow6 = (X5bow6 & E6bow6);
assign E6bow6 = (~(Ssaow6 & Evyiu6));
assign Ssaow6 = (L6bow6 & Y31ju6);
assign L6bow6 = (~(Xkaow6 | D7fpw6[15]));
assign X5bow6 = (Ax1ju6 | Ad8iu6);
assign Puaow6 = (S6bow6 & Z6bow6);
assign Z6bow6 = (G7bow6 & N7bow6);
assign N7bow6 = (~(Omyiu6 & U7bow6));
assign U7bow6 = (~(B8bow6 & I8bow6));
assign I8bow6 = (P8bow6 & W8bow6);
assign W8bow6 = (~(Apaiu6 & D9bow6));
assign D9bow6 = (~(K9bow6 & R9bow6));
assign R9bow6 = (~(Y9bow6 & Tfjiu6));
assign Y9bow6 = (Y2oiu6 | P0biu6);
assign P8bow6 = (Fabow6 & Mabow6);
assign Mabow6 = (~(Tabow6 & T4aow6));
assign T4aow6 = (Abbow6 & Hbbow6);
assign Abbow6 = (Ya1ju6 & Frziu6);
assign Tabow6 = (~(G7oiu6 | Qpaju6));
assign Fabow6 = (~(Obbow6 & Vbbow6));
assign Vbbow6 = (Wp0iu6 | Ep6ow6);
assign Ep6ow6 = (Taaiu6 & Tr0iu6);
assign B8bow6 = (Ccbow6 & Jcbow6);
assign Jcbow6 = (~(Qcbow6 & Ruaiu6));
assign Qcbow6 = (~(Xcbow6 & Edbow6));
assign Edbow6 = (~(Sy2ju6 & Kxziu6));
assign Sy2ju6 = (Cyfpw6[4] & Mr0iu6);
assign Xcbow6 = (P1bow6 | Knaiu6);
assign Ccbow6 = (~(Oxniu6 & Pugiu6));
assign Oxniu6 = (Cyfpw6[0] & Zraiu6);
assign G7bow6 = (Ax1ju6 | D7fpw6[7]);
assign Ax1ju6 = (~(Ldbow6 & Z4jiu6));
assign Z4jiu6 = (~(Hujiu6 | Gkiiu6));
assign Ldbow6 = (Htyiu6 & Sdbow6);
assign Htyiu6 = (W0piu6 & Geaiu6);
assign S6bow6 = (~(Zdbow6 | Gebow6));
assign Gebow6 = (~(R2aiu6 | Lkaiu6));
assign Zdbow6 = (Cyfpw6[7] ? Nebow6 : Mfjiu6);
assign Nebow6 = (~(Uebow6 & Bfbow6));
assign Bfbow6 = (~(D6kiu6 & Pugiu6));
assign Uebow6 = (Ifbow6 & Pfbow6);
assign Pfbow6 = (~(I82ju6 & Xojiu6));
assign Ifbow6 = (~(Jf6ju6 & It2ju6));
assign Oqohu6 = (~(Wfbow6 & Dgbow6));
assign Dgbow6 = (~(Y7ghu6 & Kgbow6));
assign Kgbow6 = (Eh6iu6 | J79ow6);
assign J79ow6 = (Ii0iu6 & Hs0iu6);
assign Wfbow6 = (~(HREADY & Rgbow6));
assign Rgbow6 = (~(Ygbow6 & Fhbow6));
assign Fhbow6 = (Mhbow6 & Thbow6);
assign Thbow6 = (Aibow6 & Hibow6);
assign Hibow6 = (~(Oibow6 & Vibow6));
assign Vibow6 = (~(D7fpw6[8] | Sbghu6));
assign Oibow6 = (Dd7ow6 & Jehhu6);
assign Dd7ow6 = (Cjbow6 & Jjbow6);
assign Jjbow6 = (J9kiu6 & D7fpw6[13]);
assign Cjbow6 = (Y40ju6 & F6ziu6);
assign Aibow6 = (~(Imaiu6 & Qjbow6));
assign Qjbow6 = (Lraiu6 | Xjbow6);
assign Mhbow6 = (Vx1ju6 & Ekbow6);
assign Ekbow6 = (~(Lkbow6 & Xe8iu6));
assign Lkbow6 = (~(Skbow6 & Zkbow6));
assign Zkbow6 = (K9aiu6 | Sbghu6);
assign Skbow6 = (Glbow6 & Nlbow6);
assign Nlbow6 = (~(Ulbow6 & Xjbow6));
assign Ulbow6 = (~(Szniu6 | Wfoiu6));
assign Szniu6 = (!Kfiiu6);
assign Kfiiu6 = (Cyfpw6[4] & K9aiu6);
assign Glbow6 = (~(Bmbow6 & E6oiu6));
assign Bmbow6 = (~(Q5aiu6 | As0iu6));
assign Vx1ju6 = (Jojiu6 | Mjfiu6);
assign Ygbow6 = (Imbow6 & Pmbow6);
assign Imbow6 = (Wmbow6 & Dnbow6);
assign Dnbow6 = (Kq0iu6 | W2aow6);
assign Wmbow6 = (Zraiu6 | Lkaiu6);
assign Hqohu6 = (F2biu6 ? B0biu6 : V9ghu6);
assign B0biu6 = (!Knbow6);
assign Aqohu6 = (G81ju6 ? H2fpw6[2] : Rnbow6);
assign Rnbow6 = (~(Ynbow6 & Fobow6));
assign Fobow6 = (Mobow6 & Tobow6);
assign Tobow6 = (~(Fb1ju6 & D7fpw6[10]));
assign Fb1ju6 = (Llaow6 & Apbow6);
assign Apbow6 = (~(Hpbow6 & Opbow6));
assign Opbow6 = (~(Vk9ow6 & D7fpw6[13]));
assign Hpbow6 = (Ftjiu6 | X1ziu6);
assign Mobow6 = (~(P91ju6 & D7fpw6[5]));
assign P91ju6 = (Llaow6 & Vpbow6);
assign Vpbow6 = (~(Cqbow6 & Jqbow6));
assign Jqbow6 = (D7fpw6[13] ? Xqbow6 : Qqbow6);
assign Xqbow6 = (~(Aujiu6 & D7fpw6[9]));
assign Qqbow6 = (Gkiiu6 | D7fpw6[15]);
assign Cqbow6 = (Erbow6 & Co6ow6);
assign Erbow6 = (Nj6ow6 | D7fpw6[12]);
assign Nj6ow6 = (D7fpw6[13] | D7fpw6[14]);
assign Ynbow6 = (Ir6ow6 & Lrbow6);
assign Lrbow6 = (~(D7fpw6[2] & Ac1ju6));
assign Ac1ju6 = (Srbow6 | Zrbow6);
assign Zrbow6 = (Gsbow6 & V4aiu6);
assign Tpohu6 = (~(Nsbow6 & Usbow6));
assign Usbow6 = (Btbow6 | Dk7ow6);
assign Nsbow6 = (Rk7ow6 ? Qjoiu6 : Itbow6);
assign Itbow6 = (Ptbow6 & Wtbow6);
assign Wtbow6 = (Dubow6 & Kubow6);
assign Kubow6 = (W6jiu6 & Faaiu6);
assign W6jiu6 = (Jc2ju6 | K9aiu6);
assign Dubow6 = (Rubow6 & Yubow6);
assign Yubow6 = (~(Fvbow6 & D7fpw6[10]));
assign Fvbow6 = (Mvbow6 & Ftjiu6);
assign Mvbow6 = (~(O8kiu6 & Tvbow6));
assign Tvbow6 = (Yb9ow6 | Qpaju6);
assign O8kiu6 = (~(Bziiu6 & Zraiu6));
assign Bziiu6 = (~(Co6ow6 | Jjhiu6));
assign Rubow6 = (~(Am7ow6 & Ppfpw6[4]));
assign Am7ow6 = (Ivfhu6 & Awbow6);
assign Awbow6 = (~(Hwbow6 & Twniu6));
assign Twniu6 = (~(D6kiu6 & Cyfpw6[1]));
assign Hwbow6 = (~(Mfjiu6 | Gsbow6));
assign Ptbow6 = (Owbow6 & Vwbow6);
assign Vwbow6 = (V4aiu6 | Cn7ow6);
assign V4aiu6 = (!D7fpw6[3]);
assign Owbow6 = (Cxbow6 & Jxbow6);
assign Jxbow6 = (A1kiu6 | Hm7ow6);
assign Cxbow6 = (~(Cbbiu6 & D7fpw6[9]));
assign Cbbiu6 = (~(Vhiiu6 | Ftjiu6));
assign Vhiiu6 = (C27ow6 | Qpaju6);
assign Mpohu6 = (~(Qxbow6 & Xxbow6));
assign Xxbow6 = (Eybow6 & Lybow6);
assign Lybow6 = (~(Egziu6 & Eafpw6[28]));
assign Eybow6 = (Sybow6 & Sgziu6);
assign Sybow6 = (Ft6ow6 | Acniu6);
assign Acniu6 = (Zybow6 & Gzbow6);
assign Gzbow6 = (Nzbow6 & Uzbow6);
assign Uzbow6 = (Iiziu6 | B0cow6);
assign Nzbow6 = (I0cow6 & Djziu6);
assign I0cow6 = (Kjziu6 | P0cow6);
assign Zybow6 = (W0cow6 & D1cow6);
assign D1cow6 = (K1cow6 | Hlziu6);
assign W0cow6 = (Mkziu6 | R1cow6);
assign Qxbow6 = (Y1cow6 & F2cow6);
assign F2cow6 = (~(Zsfpw6[27] & Cmziu6));
assign Y1cow6 = (~(vis_pc_o[27] & Jmziu6));
assign Fpohu6 = (~(M2cow6 & T2cow6));
assign T2cow6 = (A3cow6 & H3cow6);
assign H3cow6 = (~(Egziu6 & Eafpw6[30]));
assign A3cow6 = (O3cow6 & Sgziu6);
assign O3cow6 = (Ft6ow6 | D5liu6);
assign D5liu6 = (V3cow6 & C4cow6);
assign C4cow6 = (J4cow6 & Q4cow6);
assign Q4cow6 = (~(X4cow6 & Rc8ow6));
assign J4cow6 = (E5cow6 & Djziu6);
assign E5cow6 = (Mkziu6 | L5cow6);
assign V3cow6 = (S5cow6 & Z5cow6);
assign Z5cow6 = (Hlziu6 | G6cow6);
assign S5cow6 = (~(N6cow6 & Dc8ow6));
assign M2cow6 = (U6cow6 & B7cow6);
assign B7cow6 = (~(Zsfpw6[29] & Cmziu6));
assign U6cow6 = (~(vis_pc_o[29] & Jmziu6));
assign Yoohu6 = (P7cow6 ? I7cow6 : Yyfhu6);
assign P7cow6 = (~(Q08iu6 | Eh6iu6));
assign Q08iu6 = (!W7cow6);
assign Roohu6 = (~(D8cow6 & K8cow6));
assign K8cow6 = (R8cow6 & Y8cow6);
assign Y8cow6 = (~(Zsfpw6[22] & Cmziu6));
assign R8cow6 = (F9cow6 & M9cow6);
assign M9cow6 = (Ft6ow6 | Lvkiu6);
assign Lvkiu6 = (T9cow6 & Aacow6);
assign Aacow6 = (Hacow6 & Oacow6);
assign Oacow6 = (Vacow6 | Q88ow6);
assign Hacow6 = (~(Cbcow6 & V78ow6));
assign T9cow6 = (Jbcow6 & Qbcow6);
assign Qbcow6 = (~(Xbcow6 & X88ow6));
assign Jbcow6 = (H78ow6 | Eccow6);
assign F9cow6 = (~(Egziu6 & Eafpw6[23]));
assign D8cow6 = (Lccow6 & Sccow6);
assign Sccow6 = (~(vis_pc_o[22] & Jmziu6));
assign Koohu6 = (~(Zccow6 & Gdcow6));
assign Gdcow6 = (Ndcow6 & Udcow6);
assign Udcow6 = (~(Egziu6 & Eafpw6[27]));
assign Ndcow6 = (Becow6 & Sgziu6);
assign Becow6 = (~(Zgziu6 & I4liu6));
assign I4liu6 = (~(Iecow6 & Pecow6));
assign Pecow6 = (Wecow6 & Dfcow6);
assign Dfcow6 = (Iiziu6 | Kfcow6);
assign Wecow6 = (Rfcow6 & Djziu6);
assign Rfcow6 = (Kjziu6 | Yfcow6);
assign Iecow6 = (Fgcow6 & Mgcow6);
assign Mgcow6 = (Mkziu6 | Tgcow6);
assign Fgcow6 = (Ahcow6 | Hlziu6);
assign Zccow6 = (Hhcow6 & Ohcow6);
assign Ohcow6 = (~(Zsfpw6[26] & Cmziu6));
assign Hhcow6 = (~(vis_pc_o[26] & Jmziu6));
assign Doohu6 = (~(Vhcow6 & Cicow6));
assign Cicow6 = (Jicow6 & Qicow6);
assign Qicow6 = (~(Egziu6 & Eafpw6[26]));
assign Jicow6 = (Xicow6 & Sgziu6);
assign Xicow6 = (~(Zgziu6 & Q1liu6));
assign Q1liu6 = (~(Ejcow6 & Ljcow6));
assign Ljcow6 = (Sjcow6 & Zjcow6);
assign Zjcow6 = (Iiziu6 | Gkcow6);
assign Iiziu6 = (!Dc8ow6);
assign Sjcow6 = (Nkcow6 & Djziu6);
assign Nkcow6 = (Kjziu6 | Ukcow6);
assign Kjziu6 = (!Rc8ow6);
assign Ejcow6 = (Blcow6 & Ilcow6);
assign Ilcow6 = (Mkziu6 | Plcow6);
assign Blcow6 = (Hlziu6 | Wlcow6);
assign Vhcow6 = (Dmcow6 & Kmcow6);
assign Kmcow6 = (~(Zsfpw6[25] & Cmziu6));
assign Dmcow6 = (~(vis_pc_o[25] & Jmziu6));
assign Wnohu6 = (~(Rmcow6 & Ymcow6));
assign Ymcow6 = (Fncow6 & Mncow6);
assign Mncow6 = (~(Egziu6 & Eafpw6[25]));
assign Fncow6 = (Tncow6 & Sgziu6);
assign Tncow6 = (~(Zgziu6 & Osliu6));
assign Osliu6 = (~(Aocow6 & Hocow6));
assign Hocow6 = (Oocow6 & Vocow6);
assign Vocow6 = (~(Dc8ow6 & Ew6ow6));
assign Oocow6 = (Cpcow6 & Djziu6);
assign Cpcow6 = (~(Rc8ow6 & Cv6ow6));
assign Aocow6 = (Jpcow6 & Qpcow6);
assign Qpcow6 = (Mkziu6 | Xv6ow6);
assign Jpcow6 = (Ou6ow6 | Hlziu6);
assign Rmcow6 = (Xpcow6 & Eqcow6);
assign Eqcow6 = (~(Zsfpw6[24] & Cmziu6));
assign Xpcow6 = (~(vis_pc_o[24] & Jmziu6));
assign Pnohu6 = (~(Lqcow6 & Sqcow6));
assign Sqcow6 = (Zqcow6 & Grcow6);
assign Grcow6 = (~(Egziu6 & Eafpw6[24]));
assign Zqcow6 = (Nrcow6 & Sgziu6);
assign Nrcow6 = (~(Zgziu6 & Nu8iu6));
assign Nu8iu6 = (~(Urcow6 & Bscow6));
assign Bscow6 = (Iscow6 & Pscow6);
assign Pscow6 = (~(Dc8ow6 & Tdliu6));
assign Dc8ow6 = (~(Wscow6 & Dtcow6));
assign Wscow6 = (Ah3ju6 | Ktcow6);
assign Iscow6 = (Rtcow6 & Djziu6);
assign Djziu6 = (~(Ytcow6 & Fucow6));
assign Fucow6 = (~(Mucow6 & Tucow6));
assign Mucow6 = (~(Fg3ju6 & Ah3ju6));
assign Ah3ju6 = (Avcow6 | Df3ju6);
assign Rtcow6 = (~(Rc8ow6 & Jfliu6));
assign Rc8ow6 = (Hvcow6 | Ovcow6);
assign Hvcow6 = (~(Fg3ju6 | Ktcow6));
assign Urcow6 = (Vvcow6 & Cwcow6);
assign Cwcow6 = (Mkziu6 | Rcliu6);
assign Vvcow6 = (Veliu6 | Hlziu6);
assign Lqcow6 = (Jwcow6 & Qwcow6);
assign Qwcow6 = (~(Zsfpw6[23] & Cmziu6));
assign Jwcow6 = (~(vis_pc_o[23] & Jmziu6));
assign Inohu6 = (~(Xwcow6 & Excow6));
assign Excow6 = (Lxcow6 & Sxcow6);
assign Sxcow6 = (~(Zsfpw6[20] & Cmziu6));
assign Lxcow6 = (Zxcow6 & Gycow6);
assign Gycow6 = (Ft6ow6 | Tyliu6);
assign Tyliu6 = (Nycow6 & Uycow6);
assign Uycow6 = (Bzcow6 & Izcow6);
assign Izcow6 = (Tkziu6 | Vacow6);
assign Bzcow6 = (Rjziu6 | Pzcow6);
assign Nycow6 = (Wzcow6 & D0dow6);
assign D0dow6 = (Alziu6 | Eccow6);
assign Wzcow6 = (Mkziu6 | Piziu6);
assign Zxcow6 = (~(Egziu6 & Eafpw6[21]));
assign Xwcow6 = (Lccow6 & K0dow6);
assign K0dow6 = (~(vis_pc_o[20] & Jmziu6));
assign Bnohu6 = (~(R0dow6 & Y0dow6));
assign Y0dow6 = (F1dow6 & M1dow6);
assign M1dow6 = (~(Zsfpw6[19] & Cmziu6));
assign F1dow6 = (T1dow6 & A2dow6);
assign A2dow6 = (Ft6ow6 | S1miu6);
assign S1miu6 = (H2dow6 & O2dow6);
assign O2dow6 = (V2dow6 & C3dow6);
assign C3dow6 = (P0cow6 | Pzcow6);
assign V2dow6 = (K1cow6 | Eccow6);
assign H2dow6 = (J3dow6 & Q3dow6);
assign Q3dow6 = (R1cow6 | Vacow6);
assign J3dow6 = (Mkziu6 | B0cow6);
assign T1dow6 = (~(Egziu6 & Eafpw6[20]));
assign R0dow6 = (Lccow6 & X3dow6);
assign X3dow6 = (~(vis_pc_o[19] & Jmziu6));
assign Umohu6 = (~(E4dow6 & L4dow6));
assign L4dow6 = (S4dow6 & Z4dow6);
assign Z4dow6 = (~(Zsfpw6[18] & Cmziu6));
assign S4dow6 = (G5dow6 & N5dow6);
assign N5dow6 = (Ft6ow6 | R4miu6);
assign R4miu6 = (U5dow6 & B6dow6);
assign B6dow6 = (I6dow6 & P6dow6);
assign P6dow6 = (Mkziu6 | Kfcow6);
assign I6dow6 = (Tgcow6 | Vacow6);
assign U5dow6 = (W6dow6 & D7dow6);
assign D7dow6 = (Ahcow6 | Eccow6);
assign W6dow6 = (Yfcow6 | Pzcow6);
assign G5dow6 = (~(Egziu6 & Eafpw6[19]));
assign E4dow6 = (Lccow6 & K7dow6);
assign K7dow6 = (~(vis_pc_o[18] & Jmziu6));
assign Nmohu6 = (~(R7dow6 & Y7dow6));
assign Y7dow6 = (F8dow6 & M8dow6);
assign M8dow6 = (~(Zsfpw6[17] & Cmziu6));
assign F8dow6 = (T8dow6 & A9dow6);
assign A9dow6 = (Ft6ow6 | Q7miu6);
assign Q7miu6 = (H9dow6 & O9dow6);
assign O9dow6 = (V9dow6 & Cadow6);
assign Cadow6 = (Vacow6 | Plcow6);
assign V9dow6 = (Pzcow6 | Ukcow6);
assign Pzcow6 = (!Cbcow6);
assign H9dow6 = (Jadow6 & Qadow6);
assign Qadow6 = (Mkziu6 | Gkcow6);
assign Mkziu6 = (!Xbcow6);
assign Jadow6 = (Eccow6 | Wlcow6);
assign T8dow6 = (~(Egziu6 & Eafpw6[18]));
assign R7dow6 = (Lccow6 & Xadow6);
assign Xadow6 = (~(vis_pc_o[17] & Jmziu6));
assign Gmohu6 = (~(Ebdow6 & Lbdow6));
assign Lbdow6 = (Sbdow6 & Zbdow6);
assign Zbdow6 = (~(Zsfpw6[16] & Cmziu6));
assign Sbdow6 = (Gcdow6 & Ncdow6);
assign Ncdow6 = (Ft6ow6 | Pamiu6);
assign Pamiu6 = (Ucdow6 & Bddow6);
assign Bddow6 = (Iddow6 & Pddow6);
assign Pddow6 = (~(Xbcow6 & Ew6ow6));
assign Iddow6 = (Xv6ow6 | Vacow6);
assign Ucdow6 = (Wddow6 & Dedow6);
assign Dedow6 = (Ou6ow6 | Eccow6);
assign Wddow6 = (~(Cv6ow6 & Cbcow6));
assign Gcdow6 = (~(Egziu6 & Eafpw6[17]));
assign Ebdow6 = (Lccow6 & Kedow6);
assign Kedow6 = (~(vis_pc_o[16] & Jmziu6));
assign Zlohu6 = (~(Redow6 & Yedow6));
assign Yedow6 = (Ffdow6 & Mfdow6);
assign Mfdow6 = (~(Zsfpw6[15] & Cmziu6));
assign Ffdow6 = (Tfdow6 & Agdow6);
assign Agdow6 = (Ft6ow6 | Odmiu6);
assign Odmiu6 = (Hgdow6 & Ogdow6);
assign Ogdow6 = (Vgdow6 & Chdow6);
assign Chdow6 = (~(Xbcow6 & Tdliu6));
assign Vgdow6 = (Rcliu6 | Vacow6);
assign Hgdow6 = (Jhdow6 & Qhdow6);
assign Qhdow6 = (Veliu6 | Eccow6);
assign Jhdow6 = (~(Jfliu6 & Cbcow6));
assign Tfdow6 = (~(Egziu6 & Eafpw6[16]));
assign Redow6 = (Lccow6 & Xhdow6);
assign Xhdow6 = (~(vis_pc_o[15] & Jmziu6));
assign Slohu6 = (~(Eidow6 & Lidow6));
assign Lidow6 = (Sidow6 & Zidow6);
assign Zidow6 = (~(Egziu6 & Eafpw6[14]));
assign Sidow6 = (Gjdow6 & Sgziu6);
assign Gjdow6 = (~(Zgziu6 & Yimiu6));
assign Yimiu6 = (~(Njdow6 & Ujdow6));
assign Ujdow6 = (Bkdow6 & Ikdow6);
assign Ikdow6 = (L5cow6 | Pkdow6);
assign Bkdow6 = (Wkdow6 & Dldow6);
assign Wkdow6 = (G6cow6 | Kldow6);
assign Njdow6 = (Rldow6 & Yldow6);
assign Yldow6 = (~(X4cow6 & Fmdow6));
assign Rldow6 = (~(N6cow6 & Mmdow6));
assign Eidow6 = (Tmdow6 & Andow6);
assign Andow6 = (~(Zsfpw6[13] & Cmziu6));
assign Tmdow6 = (~(vis_pc_o[13] & Jmziu6));
assign Llohu6 = (~(Hndow6 & Ondow6));
assign Ondow6 = (Vndow6 & Codow6);
assign Codow6 = (~(Egziu6 & Eafpw6[13]));
assign Vndow6 = (Jodow6 & Sgziu6);
assign Jodow6 = (~(Zgziu6 & Qlmiu6));
assign Qlmiu6 = (~(Qodow6 & Xodow6));
assign Xodow6 = (Epdow6 & Lpdow6);
assign Lpdow6 = (Rjziu6 | Spdow6);
assign Epdow6 = (Zpdow6 & Dldow6);
assign Zpdow6 = (Tkziu6 | Pkdow6);
assign Qodow6 = (Gqdow6 & Nqdow6);
assign Nqdow6 = (Alziu6 | Kldow6);
assign Gqdow6 = (Piziu6 | Uqdow6);
assign Hndow6 = (Brdow6 & Irdow6);
assign Irdow6 = (~(Zsfpw6[12] & Cmziu6));
assign Brdow6 = (~(vis_pc_o[12] & Jmziu6));
assign Elohu6 = (~(Prdow6 & Wrdow6));
assign Wrdow6 = (Dsdow6 & Ksdow6);
assign Ksdow6 = (~(Egziu6 & Eafpw6[12]));
assign Dsdow6 = (Rsdow6 & Sgziu6);
assign Rsdow6 = (~(Zgziu6 & Iomiu6));
assign Iomiu6 = (~(Ysdow6 & Ftdow6));
assign Ftdow6 = (Mtdow6 & Ttdow6);
assign Ttdow6 = (K1cow6 | Kldow6);
assign Mtdow6 = (Audow6 & Dldow6);
assign Audow6 = (P0cow6 | Spdow6);
assign Ysdow6 = (Hudow6 & Oudow6);
assign Oudow6 = (R1cow6 | Pkdow6);
assign Hudow6 = (B0cow6 | Uqdow6);
assign Prdow6 = (Vudow6 & Cvdow6);
assign Cvdow6 = (~(Zsfpw6[11] & Cmziu6));
assign Vudow6 = (~(vis_pc_o[11] & Jmziu6));
assign Xkohu6 = (~(Jvdow6 & Qvdow6));
assign Qvdow6 = (Xvdow6 & Ewdow6);
assign Ewdow6 = (~(Egziu6 & Eafpw6[8]));
assign Xvdow6 = (Lwdow6 & Sgziu6);
assign Lwdow6 = (~(Zgziu6 & E7niu6));
assign E7niu6 = (~(Swdow6 & Zwdow6));
assign Zwdow6 = (Gxdow6 & Nxdow6);
assign Nxdow6 = (Rcliu6 | Pkdow6);
assign Rcliu6 = (Uxdow6 & Bydow6);
assign Bydow6 = (Iydow6 | W4siu6);
assign W4siu6 = (Pydow6 & Wydow6);
assign Wydow6 = (Dzdow6 & Kzdow6);
assign Kzdow6 = (~(Tzfpw6[8] & Yvgiu6));
assign Dzdow6 = (Rzdow6 & Yzdow6);
assign Yzdow6 = (~(F0eow6 & Vbgpw6[8]));
assign Rzdow6 = (~(M0eow6 & Odgpw6[8]));
assign Pydow6 = (T0eow6 & A1eow6);
assign A1eow6 = (~(Bagpw6[8] & M6eiu6));
assign T0eow6 = (~(STCALIB[8] & H1eow6));
assign Uxdow6 = (O1eow6 & V1eow6);
assign V1eow6 = (~(Gk3ju6 & C2eow6));
assign Gk3ju6 = (J2eow6 ? Cw3ju6 : Tf4ju6);
assign O1eow6 = (~(HRDATA[8] & Q2eow6));
assign Gxdow6 = (X2eow6 & Dldow6);
assign X2eow6 = (~(Tdliu6 & Mmdow6));
assign Tdliu6 = (~(E3eow6 & L3eow6));
assign L3eow6 = (Iydow6 | M1xiu6);
assign M1xiu6 = (S3eow6 & Z3eow6);
assign Z3eow6 = (G4eow6 & N4eow6);
assign N4eow6 = (U4eow6 & B5eow6);
assign B5eow6 = (~(STCALIB[0] & H1eow6));
assign U4eow6 = (~(ECOREVNUM[0] & I5eow6));
assign G4eow6 = (P5eow6 & W5eow6);
assign W5eow6 = (~(Y5eiu6 & Bxghu6));
assign P5eow6 = (~(Yvgiu6 & Tzfpw6[0]));
assign S3eow6 = (D6eow6 & K6eow6);
assign K6eow6 = (R6eow6 & Y6eow6);
assign Y6eow6 = (~(Bagpw6[0] & M6eiu6));
assign R6eow6 = (~(Odgpw6[0] & M0eow6));
assign D6eow6 = (F7eow6 & M7eow6);
assign M7eow6 = (~(T7eow6 & vis_ipsr_o[0]));
assign F7eow6 = (~(F0eow6 & Vbgpw6[0]));
assign E3eow6 = (A8eow6 & H8eow6);
assign H8eow6 = (~(C2eow6 & Lj3ju6));
assign Lj3ju6 = (Hv3ju6 ? Sx3ju6 : O8eow6);
assign A8eow6 = (~(HRDATA[0] & Q2eow6));
assign Swdow6 = (V8eow6 & C9eow6);
assign C9eow6 = (Veliu6 | Kldow6);
assign Veliu6 = (J9eow6 & Q9eow6);
assign Q9eow6 = (Iydow6 | Gntiu6);
assign Gntiu6 = (X9eow6 & Eaeow6);
assign Eaeow6 = (Laeow6 & Saeow6);
assign Saeow6 = (Zaeow6 & Gbeow6);
assign Gbeow6 = (~(Bagpw6[16] & M6eiu6));
assign Zaeow6 = (~(Tzfpw6[16] & Yvgiu6));
assign Laeow6 = (Nbeow6 & Ubeow6);
assign Ubeow6 = (~(Krghu6 & Y5eiu6));
assign Nbeow6 = (~(Odgpw6[16] & M0eow6));
assign X9eow6 = (Bceow6 & Iceow6);
assign Iceow6 = (~(Pceow6 & Wceow6));
assign Wceow6 = (Nzhiu6 | Vbgpw6[16]);
assign Bceow6 = (Ddeow6 & Kdeow6);
assign Kdeow6 = (~(STCALIB[16] & H1eow6));
assign Ddeow6 = (Z4ciu6 | Qkgiu6);
assign Z4ciu6 = (~(Rdeow6 & Ydeow6));
assign Rdeow6 = (~(Feeow6 | Meeow6));
assign J9eow6 = (Teeow6 & Afeow6);
assign Afeow6 = (Uk3ju6 | Hfeow6);
assign Uk3ju6 = (!Ofeow6);
assign Ofeow6 = (Hv3ju6 ? E44ju6 : Ke4ju6);
assign Teeow6 = (~(HRDATA[16] & Q2eow6));
assign V8eow6 = (~(Jfliu6 & Fmdow6));
assign Jfliu6 = (~(Vfeow6 & Cgeow6));
assign Cgeow6 = (Iydow6 | P8viu6);
assign P8viu6 = (Jgeow6 & Qgeow6);
assign Jgeow6 = (Xgeow6 & Eheow6);
assign Eheow6 = (~(M0eow6 & Odgpw6[24]));
assign Xgeow6 = (~(F0eow6 & Vbgpw6[24]));
assign Vfeow6 = (Lheow6 & Sheow6);
assign Sheow6 = (~(HRDATA[24] & Q2eow6));
assign Lheow6 = (~(C2eow6 & Eb4ju6));
assign Eb4ju6 = (~(Zheow6 & Gieow6));
assign Gieow6 = (~(Nieow6 & Vh3ju6));
assign Zheow6 = (Nk3ju6 | Nieow6);
assign Nieow6 = (~(Uieow6 | Ii0iu6));
assign Nk3ju6 = (!Bjeow6);
assign Bjeow6 = (Hv3ju6 ? Ijeow6 : V24ju6);
assign Jvdow6 = (Pjeow6 & Wjeow6);
assign Wjeow6 = (~(Zsfpw6[7] & Cmziu6));
assign Pjeow6 = (~(vis_pc_o[7] & Jmziu6));
assign Qkohu6 = (~(Dkeow6 & Kkeow6));
assign Kkeow6 = (Rkeow6 & Ykeow6);
assign Ykeow6 = (~(Egziu6 & Eafpw6[6]));
assign Rkeow6 = (Fleow6 & Sgziu6);
assign Fleow6 = (~(Zgziu6 & Wqkiu6));
assign Wqkiu6 = (~(Mleow6 & Tleow6));
assign Tleow6 = (Ameow6 & Hmeow6);
assign Hmeow6 = (Cfliu6 | G6cow6);
assign Ameow6 = (Omeow6 & Mdliu6);
assign Omeow6 = (~(Qfliu6 & X4cow6));
assign Mleow6 = (Vmeow6 & Cneow6);
assign Cneow6 = (Ycliu6 | L5cow6);
assign Vmeow6 = (~(Aeliu6 & N6cow6));
assign Dkeow6 = (Jneow6 & Qneow6);
assign Qneow6 = (~(Zsfpw6[5] & Cmziu6));
assign Jneow6 = (~(vis_pc_o[5] & Jmziu6));
assign Jkohu6 = (~(Xneow6 & Eoeow6));
assign Eoeow6 = (Loeow6 & Soeow6);
assign Soeow6 = (~(Egziu6 & Eafpw6[5]));
assign Loeow6 = (Zoeow6 & Sgziu6);
assign Zoeow6 = (Ft6ow6 | Ljbiu6);
assign Ljbiu6 = (Gpeow6 & Npeow6);
assign Npeow6 = (Upeow6 & Bqeow6);
assign Bqeow6 = (Rjziu6 | Iqeow6);
assign Rjziu6 = (Pqeow6 & Wqeow6);
assign Wqeow6 = (Iydow6 | U6wiu6);
assign U6wiu6 = (Dreow6 & Kreow6);
assign Kreow6 = (~(F0eow6 & Vbgpw6[29]));
assign Dreow6 = (Rreow6 & Yreow6);
assign Rreow6 = (~(Odgpw6[29] & M0eow6));
assign Pqeow6 = (Fseow6 & Mseow6);
assign Mseow6 = (~(C2eow6 & Tseow6));
assign Tseow6 = (~(T84ju6 & Ateow6));
assign Ateow6 = (Hteow6 | Bz3ju6);
assign T84ju6 = (~(Oteow6 & Vteow6));
assign Vteow6 = (Ex3ju6 | J2eow6);
assign Oteow6 = (Cueow6 & Hteow6);
assign Hteow6 = (~(Jueow6 & Queow6));
assign Jueow6 = (Xueow6 & Eveow6);
assign Eveow6 = (~(Lveow6 & Sveow6));
assign Xueow6 = (Zveow6 | Gweow6);
assign Cueow6 = (~(Nweow6 & J2eow6));
assign Fseow6 = (~(Q2eow6 & HRDATA[29]));
assign Upeow6 = (Uweow6 & Mdliu6);
assign Uweow6 = (Tkziu6 | Ycliu6);
assign Tkziu6 = (Bxeow6 & Ixeow6);
assign Ixeow6 = (Pxeow6 & Wxeow6);
assign Wxeow6 = (~(Dyeow6 & Ff4ju6));
assign Pxeow6 = (Iydow6 | U2tiu6);
assign U2tiu6 = (Kyeow6 & Ryeow6);
assign Ryeow6 = (Yyeow6 & Fzeow6);
assign Fzeow6 = (~(Tzfpw6[13] & Yvgiu6));
assign Yyeow6 = (Mzeow6 & Tzeow6);
assign Tzeow6 = (~(T7eow6 & E4ciu6));
assign E4ciu6 = (~(A0fow6 & H0fow6));
assign H0fow6 = (~(O0fow6 & V0fow6));
assign O0fow6 = (~(C1fow6 & J1fow6));
assign C1fow6 = (E2fow6 ? X1fow6 : Q1fow6);
assign X1fow6 = (L2fow6 & S2fow6);
assign S2fow6 = (~(Z2fow6 & G3fow6));
assign L2fow6 = (B4fow6 ? U3fow6 : N3fow6);
assign U3fow6 = (I4fow6 | P4fow6);
assign N3fow6 = (K5fow6 ? D5fow6 : W4fow6);
assign Q1fow6 = (R5fow6 & Y5fow6);
assign Y5fow6 = (F6fow6 | M6fow6);
assign R5fow6 = (H7fow6 ? A7fow6 : T6fow6);
assign A7fow6 = (O7fow6 | V7fow6);
assign T6fow6 = (~(C8fow6 | J8fow6));
assign J8fow6 = (~(Q8fow6 | X8fow6));
assign Mzeow6 = (~(Odgpw6[13] & M0eow6));
assign Kyeow6 = (E9fow6 & L9fow6);
assign L9fow6 = (~(F0eow6 & Vbgpw6[13]));
assign E9fow6 = (S9fow6 & Z9fow6);
assign Z9fow6 = (~(STCALIB[13] & H1eow6));
assign S9fow6 = (~(Bagpw6[13] & M6eiu6));
assign Bxeow6 = (Gafow6 & Nafow6);
assign Nafow6 = (Uafow6 | Uc4ju6);
assign Gafow6 = (~(Q2eow6 & HRDATA[13]));
assign Gpeow6 = (Bbfow6 & Ibfow6);
assign Ibfow6 = (Alziu6 | Cfliu6);
assign Alziu6 = (Pbfow6 & Wbfow6);
assign Wbfow6 = (Dcfow6 & Kcfow6);
assign Kcfow6 = (Rcfow6 | J34ju6);
assign J34ju6 = (!V94ju6);
assign Dcfow6 = (Iydow6 | Umuiu6);
assign Umuiu6 = (Ycfow6 & Fdfow6);
assign Fdfow6 = (Mdfow6 & Tdfow6);
assign Tdfow6 = (~(Tzfpw6[21] & Yvgiu6));
assign Mdfow6 = (Aefow6 & Hefow6);
assign Hefow6 = (~(F0eow6 & Vbgpw6[21]));
assign Aefow6 = (~(Odgpw6[21] & M0eow6));
assign Ycfow6 = (Oefow6 & Vefow6);
assign Vefow6 = (~(Bagpw6[21] & M6eiu6));
assign Oefow6 = (~(STCALIB[21] & H1eow6));
assign Pbfow6 = (Cffow6 & Jffow6);
assign Jffow6 = (Uafow6 | F14ju6);
assign Cffow6 = (~(HRDATA[21] & Q2eow6));
assign Bbfow6 = (Piziu6 | Qffow6);
assign Piziu6 = (Xffow6 & Egfow6);
assign Egfow6 = (Lgfow6 & Sgfow6);
assign Sgfow6 = (~(Dyeow6 & Hg4ju6));
assign Lgfow6 = (Iydow6 | Eariu6);
assign Eariu6 = (Zgfow6 & Ghfow6);
assign Ghfow6 = (Nhfow6 & Uhfow6);
assign Uhfow6 = (~(Tzfpw6[5] & Yvgiu6));
assign Nhfow6 = (Bifow6 & Iifow6);
assign Iifow6 = (~(Bagpw6[5] & M6eiu6));
assign Bifow6 = (~(Odgpw6[5] & M0eow6));
assign Zgfow6 = (Pifow6 & Wifow6);
assign Wifow6 = (~(F0eow6 & Vbgpw6[5]));
assign Pifow6 = (Djfow6 & Kjfow6);
assign Kjfow6 = (~(STCALIB[5] & H1eow6));
assign Djfow6 = (Qkgiu6 | Vhbiu6);
assign Xffow6 = (Rjfow6 & Yjfow6);
assign Yjfow6 = (Uafow6 | Mu3ju6);
assign Rjfow6 = (~(HRDATA[5] & Q2eow6));
assign Xneow6 = (Fkfow6 & Mkfow6);
assign Mkfow6 = (~(Zsfpw6[4] & Cmziu6));
assign Fkfow6 = (~(vis_pc_o[4] & Jmziu6));
assign Ckohu6 = (~(Tkfow6 & Alfow6));
assign Alfow6 = (Hlfow6 & Olfow6);
assign Olfow6 = (~(Egziu6 & Eafpw6[4]));
assign Hlfow6 = (Vlfow6 & Sgziu6);
assign Vlfow6 = (Ft6ow6 | Y4fiu6);
assign Y4fiu6 = (Cmfow6 & Jmfow6);
assign Jmfow6 = (Qmfow6 & Xmfow6);
assign Xmfow6 = (K1cow6 | Cfliu6);
assign K1cow6 = (Enfow6 & Lnfow6);
assign Lnfow6 = (Snfow6 & Znfow6);
assign Znfow6 = (~(Dyeow6 & V24ju6));
assign V24ju6 = (~(Gofow6 & Nofow6));
assign Nofow6 = (Uofow6 & Bpfow6);
assign Bpfow6 = (Ipfow6 | A70iu6);
assign Uofow6 = (Ppfow6 | V70iu6);
assign Gofow6 = (Wpfow6 & Dqfow6);
assign Dqfow6 = (Kqfow6 | O70iu6);
assign Wpfow6 = (Rqfow6 | H70iu6);
assign Snfow6 = (Iydow6 | Bguiu6);
assign Bguiu6 = (Yqfow6 & Frfow6);
assign Frfow6 = (Mrfow6 & Trfow6);
assign Trfow6 = (~(Tzfpw6[20] & Yvgiu6));
assign Mrfow6 = (Asfow6 & Hsfow6);
assign Hsfow6 = (~(F0eow6 & Vbgpw6[20]));
assign Asfow6 = (~(Odgpw6[20] & M0eow6));
assign Yqfow6 = (Osfow6 & Vsfow6);
assign Vsfow6 = (~(Bagpw6[20] & M6eiu6));
assign Osfow6 = (~(STCALIB[20] & H1eow6));
assign Enfow6 = (Ctfow6 & Jtfow6);
assign Jtfow6 = (~(Qtfow6 & E44ju6));
assign E44ju6 = (~(Xtfow6 & Eufow6));
assign Eufow6 = (Lufow6 & Sufow6);
assign Sufow6 = (Ipfow6 | C80iu6);
assign Lufow6 = (Rqfow6 | J80iu6);
assign Xtfow6 = (Zufow6 & Gvfow6);
assign Gvfow6 = (Ppfow6 | X80iu6);
assign Zufow6 = (Kqfow6 | Q80iu6);
assign Ctfow6 = (~(HRDATA[20] & Q2eow6));
assign Qmfow6 = (Nvfow6 & Mdliu6);
assign Nvfow6 = (P0cow6 | Iqeow6);
assign P0cow6 = (Uvfow6 & Bwfow6);
assign Bwfow6 = (Iydow6 | I0wiu6);
assign I0wiu6 = (Iwfow6 & Pwfow6);
assign Pwfow6 = (~(Pceow6 & Wwfow6));
assign Wwfow6 = (Nzhiu6 | Vbgpw6[28]);
assign Iwfow6 = (Dxfow6 & Kxfow6);
assign Kxfow6 = (Jh5iu6 | Qkgiu6);
assign Jh5iu6 = (!Ikghu6);
assign Dxfow6 = (~(Odgpw6[28] & M0eow6));
assign Uvfow6 = (Rxfow6 & Yxfow6);
assign Yxfow6 = (~(C2eow6 & Xa4ju6));
assign Xa4ju6 = (Myfow6 ? Vh3ju6 : Fyfow6);
assign Myfow6 = (Tyfow6 & Cyfpw6[3]);
assign Tyfow6 = (Azfow6 & Hzfow6);
assign Fyfow6 = (Hv3ju6 ? O8eow6 : Ijeow6);
assign O8eow6 = (~(Ozfow6 & Vzfow6));
assign Vzfow6 = (C0gow6 & J0gow6);
assign J0gow6 = (Rqfow6 | F60iu6);
assign C0gow6 = (Ipfow6 | K50iu6);
assign Ozfow6 = (Q0gow6 & X0gow6);
assign X0gow6 = (Ppfow6 | Dc0iu6);
assign Q0gow6 = (Kqfow6 | E90iu6);
assign Ijeow6 = (~(E1gow6 & L1gow6));
assign L1gow6 = (S1gow6 & Z1gow6);
assign Z1gow6 = (Ipfow6 | R50iu6);
assign S1gow6 = (Ppfow6 | T60iu6);
assign E1gow6 = (G2gow6 & N2gow6);
assign N2gow6 = (Kqfow6 | M60iu6);
assign G2gow6 = (Rqfow6 | Y50iu6);
assign Rxfow6 = (~(HRDATA[28] & Q2eow6));
assign Cmfow6 = (U2gow6 & B3gow6);
assign B3gow6 = (R1cow6 | Ycliu6);
assign R1cow6 = (I3gow6 & P3gow6);
assign P3gow6 = (W3gow6 & D4gow6);
assign D4gow6 = (~(Dyeow6 & Ke4ju6));
assign Ke4ju6 = (~(K4gow6 & R4gow6));
assign R4gow6 = (Y4gow6 & F5gow6);
assign F5gow6 = (Ipfow6 | L90iu6);
assign Y4gow6 = (Rqfow6 | S90iu6);
assign K4gow6 = (M5gow6 & T5gow6);
assign T5gow6 = (Ppfow6 | Ga0iu6);
assign M5gow6 = (Kqfow6 | Z90iu6);
assign W3gow6 = (Iydow6 | Nvsiu6);
assign Nvsiu6 = (A6gow6 & H6gow6);
assign H6gow6 = (O6gow6 & V6gow6);
assign V6gow6 = (~(Bagpw6[12] & M6eiu6));
assign O6gow6 = (C7gow6 & J7gow6);
assign J7gow6 = (Kmbiu6 | Qkgiu6);
assign Kmbiu6 = (~(Q7gow6 & Te6iu6));
assign Q7gow6 = (~(X7gow6 & E8gow6));
assign E8gow6 = (~(L8gow6 & S8gow6));
assign S8gow6 = (Z8gow6 | Feeow6);
assign Z8gow6 = (Meeow6 ? N9gow6 : G9gow6);
assign N9gow6 = (H7fow6 ? Bagow6 : U9gow6);
assign Bagow6 = (O7fow6 ? Pagow6 : Iagow6);
assign Pagow6 = (M6fow6 ? Dbgow6 : Wagow6);
assign Iagow6 = (V7fow6 ? Rbgow6 : Kbgow6);
assign U9gow6 = (~(Ybgow6 & Fcgow6));
assign Fcgow6 = (~(C8fow6 & Mcgow6));
assign Ybgow6 = (Hdgow6 ? Adgow6 : Tcgow6);
assign Adgow6 = (Cegow6 ? Vdgow6 : Odgow6);
assign Tcgow6 = (Jegow6 | Qegow6);
assign G9gow6 = (!Xegow6);
assign Xegow6 = (Sfgow6 ? Lfgow6 : Efgow6);
assign Lfgow6 = (Nggow6 ? Gggow6 : Zfgow6);
assign Gggow6 = (Ihgow6 ? Bhgow6 : Uggow6);
assign Zfgow6 = (Digow6 ? Whgow6 : Phgow6);
assign Efgow6 = (Yigow6 ? Rigow6 : Kigow6);
assign Rigow6 = (Tjgow6 ? Mjgow6 : Fjgow6);
assign Kigow6 = (G3fow6 ? Hkgow6 : Akgow6);
assign L8gow6 = (Okgow6 & V0fow6);
assign C7gow6 = (~(Tzfpw6[12] & Yvgiu6));
assign A6gow6 = (Vkgow6 & Clgow6);
assign Clgow6 = (~(F0eow6 & Vbgpw6[12]));
assign Vkgow6 = (Jlgow6 & Qlgow6);
assign Qlgow6 = (~(STCALIB[12] & H1eow6));
assign Jlgow6 = (~(Odgpw6[12] & M0eow6));
assign I3gow6 = (Xlgow6 & Emgow6);
assign Emgow6 = (~(Qtfow6 & Tf4ju6));
assign Tf4ju6 = (~(Lmgow6 & Smgow6));
assign Smgow6 = (Zmgow6 & Gngow6);
assign Gngow6 = (Ipfow6 | Na0iu6);
assign Zmgow6 = (Rqfow6 | Ua0iu6);
assign Lmgow6 = (Nngow6 & Ungow6);
assign Ungow6 = (Ppfow6 | Ib0iu6);
assign Nngow6 = (Kqfow6 | Bb0iu6);
assign Xlgow6 = (~(HRDATA[12] & Q2eow6));
assign U2gow6 = (B0cow6 | Qffow6);
assign B0cow6 = (Bogow6 & Iogow6);
assign Iogow6 = (Pogow6 & Wogow6);
assign Wogow6 = (~(Dyeow6 & Cw3ju6));
assign Cw3ju6 = (~(Dpgow6 & Kpgow6));
assign Kpgow6 = (Rpgow6 & Ypgow6);
assign Ypgow6 = (Ppfow6 | B40iu6);
assign Rpgow6 = (Ipfow6 | Pb0iu6);
assign Dpgow6 = (Fqgow6 & Mqgow6);
assign Mqgow6 = (Rqfow6 | Wb0iu6);
assign Fqgow6 = (Kqfow6 | U30iu6);
assign Pogow6 = (Iydow6 | Yzqiu6);
assign Yzqiu6 = (Tqgow6 & Argow6);
assign Argow6 = (Hrgow6 & Orgow6);
assign Orgow6 = (Vrgow6 & Csgow6);
assign Csgow6 = (~(Odgpw6[4] & M0eow6));
assign Vrgow6 = (~(STCALIB[4] & H1eow6));
assign Hrgow6 = (Jsgow6 & Qsgow6);
assign Qsgow6 = (~(T7eow6 & vis_ipsr_o[4]));
assign Jsgow6 = (~(F0eow6 & Vbgpw6[4]));
assign Tqgow6 = (Xsgow6 & Etgow6);
assign Etgow6 = (~(Fpgiu6 & Gfghu6));
assign Xsgow6 = (Ltgow6 & Stgow6);
assign Stgow6 = (~(Bagpw6[4] & M6eiu6));
assign Ltgow6 = (~(Tzfpw6[4] & Yvgiu6));
assign Bogow6 = (Ztgow6 & Gugow6);
assign Gugow6 = (~(Qtfow6 & Sx3ju6));
assign Sx3ju6 = (~(Nugow6 & Uugow6));
assign Uugow6 = (Bvgow6 & Ivgow6);
assign Ivgow6 = (Ipfow6 | I40iu6);
assign Bvgow6 = (Kqfow6 | W40iu6);
assign Nugow6 = (Pvgow6 & Wvgow6);
assign Wvgow6 = (Ppfow6 | D50iu6);
assign Pvgow6 = (Rqfow6 | P40iu6);
assign Ztgow6 = (~(HRDATA[4] & Q2eow6));
assign Tkfow6 = (Dwgow6 & Kwgow6);
assign Kwgow6 = (~(Zsfpw6[3] & Cmziu6));
assign Dwgow6 = (~(vis_pc_o[3] & Jmziu6));
assign Vjohu6 = (~(Rwgow6 & Ywgow6));
assign Ywgow6 = (Fxgow6 & Mxgow6);
assign Mxgow6 = (~(Egziu6 & Eafpw6[3]));
assign Fxgow6 = (Txgow6 & Sgziu6);
assign Txgow6 = (Ft6ow6 | Kifiu6);
assign Kifiu6 = (Aygow6 & Hygow6);
assign Hygow6 = (Oygow6 & Vygow6);
assign Vygow6 = (Cfliu6 | Ahcow6);
assign Oygow6 = (Czgow6 & Mdliu6);
assign Czgow6 = (Iqeow6 | Yfcow6);
assign Aygow6 = (Jzgow6 & Qzgow6);
assign Qzgow6 = (Ycliu6 | Tgcow6);
assign Jzgow6 = (Qffow6 | Kfcow6);
assign Rwgow6 = (Xzgow6 & E0how6);
assign E0how6 = (~(Zsfpw6[2] & Cmziu6));
assign Xzgow6 = (~(vis_pc_o[2] & Jmziu6));
assign Ojohu6 = (~(L0how6 & S0how6));
assign S0how6 = (Z0how6 & G1how6);
assign G1how6 = (~(Egziu6 & Eafpw6[2]));
assign Z0how6 = (N1how6 & Sgziu6);
assign N1how6 = (Ft6ow6 | Ogciu6);
assign Ogciu6 = (U1how6 & B2how6);
assign B2how6 = (I2how6 & P2how6);
assign P2how6 = (Cfliu6 | Wlcow6);
assign Cfliu6 = (W2how6 & D3how6);
assign D3how6 = (K3how6 | R3how6);
assign W2how6 = (Y3how6 & F4how6);
assign Y3how6 = (~(M4how6 & T4how6));
assign M4how6 = (~(Iwfpw6[0] | Y7ghu6));
assign I2how6 = (A5how6 & Mdliu6);
assign Mdliu6 = (~(H5how6 & O5how6));
assign O5how6 = (~(V5how6 & C6how6));
assign V5how6 = (~(J6how6 & Q6how6));
assign Q6how6 = (Ny3ju6 & Tucow6);
assign J6how6 = (Z44ju6 & X6how6);
assign Z44ju6 = (R3how6 | E7how6);
assign E7how6 = (Avcow6 & L7how6);
assign A5how6 = (Iqeow6 | Ukcow6);
assign Iqeow6 = (!Qfliu6);
assign Qfliu6 = (~(S7how6 & Z7how6));
assign Z7how6 = (~(G8how6 & Iwfpw6[1]));
assign S7how6 = (N8how6 & Dtcow6);
assign N8how6 = (X6how6 | Ktcow6);
assign U1how6 = (U8how6 & B9how6);
assign B9how6 = (Ycliu6 | Plcow6);
assign Ycliu6 = (I9how6 & P9how6);
assign P9how6 = (W9how6 & Dahow6);
assign I9how6 = (Kahow6 & Rahow6);
assign Kahow6 = (~(G8how6 & Yahow6));
assign G8how6 = (Fbhow6 & Mbhow6);
assign Mbhow6 = (~(Cyfpw6[1] | Y7ghu6));
assign Fbhow6 = (~(Tbhow6 | Tucow6));
assign Tbhow6 = (!Iwfpw6[0]);
assign U8how6 = (Qffow6 | Gkcow6);
assign Qffow6 = (!Aeliu6);
assign Aeliu6 = (~(Eccow6 & Achow6));
assign Achow6 = (~(Ktcow6 & Hchow6));
assign Hchow6 = (~(Ochow6 & Vchow6));
assign Vchow6 = (Cdhow6 & Eu0iu6);
assign Eu0iu6 = (!Jdhow6);
assign Cdhow6 = (~(Qdhow6 & Xdhow6));
assign Xdhow6 = (~(Cyfpw6[1] & Eehow6));
assign Eehow6 = (Cyfpw6[0] | Cyfpw6[3]);
assign Qdhow6 = (~(Iwfpw6[0] | Iwfpw6[1]));
assign Ochow6 = (Cyfpw6[5] & Lehow6);
assign Lehow6 = (Nlaiu6 | Tfjiu6);
assign L0how6 = (Sehow6 & Zehow6);
assign Zehow6 = (~(Zsfpw6[1] & Cmziu6));
assign Sehow6 = (Quzhu6 | Ar8iu6);
assign Quzhu6 = (!vis_pc_o[1]);
assign Hjohu6 = (~(Gfhow6 & Nfhow6));
assign Nfhow6 = (~(Ufhow6 & Ophiu6));
assign Ufhow6 = (~(Juzhu6 & Bghow6));
assign Bghow6 = (N6piu6 | Eh6iu6);
assign Gfhow6 = (~(Sufpw6[1] & Eh6iu6));
assign Ajohu6 = (!Ighow6);
assign Ighow6 = (F2biu6 ? X5phu6 : Sijiu6);
assign F2biu6 = (~(Eh6iu6 | K9aiu6));
assign X5phu6 = (~(Ivfhu6 & Pghow6));
assign Pghow6 = (~(Wghow6 & Dhhow6));
assign Dhhow6 = (Khhow6 & Rhhow6);
assign Rhhow6 = (~(Ppfpw6[8] | Ppfpw6[9]));
assign Khhow6 = (~(Ppfpw6[6] | Ppfpw6[7]));
assign Wghow6 = (Yhhow6 & Fihow6);
assign Fihow6 = (~(Ppfpw6[12] | Ppfpw6[13]));
assign Yhhow6 = (~(Ppfpw6[10] | Ppfpw6[11]));
assign Tiohu6 = (Eh6iu6 ? T6ehu6 : Mihow6);
assign Mihow6 = (~(Tihow6 & Ajhow6));
assign Ajhow6 = (~(H4oiu6 & Hjhow6));
assign Hjhow6 = (~(Xkaow6 | R75iu6));
assign H4oiu6 = (~(K9bow6 | G7oiu6));
assign Tihow6 = (~(Ojhow6 & Vjhow6));
assign Ojhow6 = (~(P1bow6 | Y2oiu6));
assign Miohu6 = (Ckhow6 | Jkhow6);
assign Jkhow6 = (~(Qkhow6 | Dk7ow6));
assign Qkhow6 = (!Xkhow6);
assign Ckhow6 = (Rk7ow6 ? S8fpw6[7] : Elhow6);
assign Elhow6 = (~(Llhow6 & Slhow6));
assign Slhow6 = (~(D7fpw6[7] & Zlhow6));
assign Llhow6 = (Ad8iu6 | Cn7ow6);
assign Fiohu6 = (Eh6iu6 ? Dxfhu6 : W7cow6);
assign Yhohu6 = (Qqhiu6 ? Hrfpw6[16] : Wz4iu6);
assign Rhohu6 = (~(Gmhow6 & Nmhow6));
assign Nmhow6 = (~(Umhow6 & HRDATA[16]));
assign Gmhow6 = (~(Hrfpw6[0] & Qqhiu6));
assign Khohu6 = (~(Bnhow6 & Inhow6));
assign Inhow6 = (~(Umhow6 & HRDATA[31]));
assign Bnhow6 = (~(Hrfpw6[15] & Qqhiu6));
assign Dhohu6 = (~(Pnhow6 & Wnhow6));
assign Wnhow6 = (~(Umhow6 & HRDATA[29]));
assign Pnhow6 = (~(Hrfpw6[13] & Qqhiu6));
assign Wgohu6 = (~(Dohow6 & Kohow6));
assign Kohow6 = (~(Umhow6 & HRDATA[28]));
assign Dohow6 = (~(Hrfpw6[12] & Qqhiu6));
assign Pgohu6 = (~(Rohow6 & Yohow6));
assign Yohow6 = (~(Umhow6 & HRDATA[27]));
assign Rohow6 = (~(Hrfpw6[11] & Qqhiu6));
assign Igohu6 = (~(Fphow6 & Mphow6));
assign Mphow6 = (~(Umhow6 & HRDATA[26]));
assign Fphow6 = (~(Hrfpw6[10] & Qqhiu6));
assign Bgohu6 = (~(Tphow6 & Aqhow6));
assign Aqhow6 = (~(Umhow6 & HRDATA[25]));
assign Tphow6 = (~(Hrfpw6[9] & Qqhiu6));
assign Ufohu6 = (~(Hqhow6 & Oqhow6));
assign Oqhow6 = (~(Umhow6 & HRDATA[24]));
assign Hqhow6 = (~(Hrfpw6[8] & Qqhiu6));
assign Nfohu6 = (~(Vqhow6 & Crhow6));
assign Crhow6 = (~(Umhow6 & HRDATA[23]));
assign Vqhow6 = (~(Hrfpw6[7] & Qqhiu6));
assign Gfohu6 = (G81ju6 ? H2fpw6[3] : Jrhow6);
assign G81ju6 = (~(HREADY & Qrhow6));
assign Qrhow6 = (~(Xrhow6 & Eshow6));
assign Eshow6 = (Lshow6 & Sshow6);
assign Sshow6 = (Zshow6 & Gthow6);
assign Gthow6 = (~(Nthow6 & Lraiu6));
assign Nthow6 = (Uu9ow6 & Uthow6);
assign Uthow6 = (~(D7fpw6[15] & Buhow6));
assign Buhow6 = (~(Iuhow6 & Bkjiu6));
assign Iuhow6 = (Rg2ju6 | D7fpw6[3]);
assign Uu9ow6 = (!X5aiu6);
assign X5aiu6 = (Puhow6 | Ttciu6);
assign Ttciu6 = (!T0hhu6);
assign Puhow6 = (E45iu6 | Ii0iu6);
assign E45iu6 = (!N20ju6);
assign Zshow6 = (~(Wuhow6 & Vviiu6));
assign Wuhow6 = (~(D7fpw6[10] | D7fpw6[8]));
assign Lshow6 = (Dvhow6 & Kvhow6);
assign Kvhow6 = (~(Y31ju6 & Rvhow6));
assign Rvhow6 = (~(Yvhow6 & Fwhow6));
assign Fwhow6 = (Mwhow6 & Twhow6);
assign Twhow6 = (~(Axhow6 & Ftjiu6));
assign Axhow6 = (~(N38ow6 & Hxhow6));
assign Hxhow6 = (~(C0ehu6 & An6ow6));
assign An6ow6 = (D7fpw6[11] | D7fpw6[7]);
assign Mwhow6 = (~(Oxhow6 | Evyiu6));
assign Oxhow6 = (Quyiu6 & Ejiiu6);
assign Ejiiu6 = (C0ehu6 & D7fpw6[12]);
assign Quyiu6 = (~(X1ziu6 | D7fpw6[11]));
assign Yvhow6 = (Vxhow6 & Cyhow6);
assign Cyhow6 = (S80ju6 | D7fpw6[8]);
assign S80ju6 = (!P0piu6);
assign Vxhow6 = (Yb9ow6 | Qxoiu6);
assign Yb9ow6 = (!Nbkiu6);
assign Dvhow6 = (~(P0piu6 & W0piu6));
assign Xrhow6 = (Jyhow6 & M1jiu6);
assign M1jiu6 = (Qyhow6 & Xyhow6);
assign Xyhow6 = (~(Ezhow6 | Wkjiu6));
assign Wkjiu6 = (Lzhow6 & Y31ju6);
assign Qyhow6 = (Szhow6 & Zzhow6);
assign Zzhow6 = (~(Hviiu6 & G0iow6));
assign G0iow6 = (~(O7ziu6 & Zt9ow6));
assign Zt9ow6 = (Od0ju6 | L01ju6);
assign Od0ju6 = (!Sdbow6);
assign Sdbow6 = (Jwiiu6 & Ndiiu6);
assign Ndiiu6 = (!D7fpw6[8]);
assign Jwiiu6 = (D7fpw6[9] & I6jiu6);
assign O7ziu6 = (!Db0ju6);
assign Szhow6 = (~(Wliiu6 & W0piu6));
assign Jyhow6 = (Onjiu6 & N0iow6);
assign N0iow6 = (Jojiu6 | Cyfpw6[7]);
assign Onjiu6 = (Yn2ju6 | Kq0iu6);
assign Jrhow6 = (~(Ir6ow6 & U0iow6));
assign U0iow6 = (~(D7fpw6[7] & B1iow6));
assign B1iow6 = (~(Uvziu6 & I1iow6));
assign I1iow6 = (~(Srbow6 & D7fpw6[10]));
assign Ir6ow6 = (P1iow6 & W1iow6);
assign W1iow6 = (D2iow6 & K2iow6);
assign K2iow6 = (~(Y7ghu6 & R2iow6));
assign R2iow6 = (Ii0iu6 | D7fpw6[3]);
assign D2iow6 = (Y2iow6 & Faaiu6);
assign Y2iow6 = (~(Aujiu6 & F3iow6));
assign F3iow6 = (Tniiu6 | Gaziu6);
assign P1iow6 = (Mb1ju6 & M3iow6);
assign M3iow6 = (~(D7fpw6[13] & Ya1ju6));
assign Mb1ju6 = (T3iow6 & A4iow6);
assign A4iow6 = (Bkjiu6 | Uvziu6);
assign Bkjiu6 = (~(R9aiu6 & D7fpw6[3]));
assign T3iow6 = (~(H4iow6 | Hs8ow6));
assign Hs8ow6 = (O4iow6 & Aujiu6);
assign O4iow6 = (~(X1ziu6 | Jcaiu6));
assign H4iow6 = (Srbow6 & V4iow6);
assign V4iow6 = (D7fpw6[11] | Q6aow6);
assign Srbow6 = (C5iow6 & J5iow6);
assign C5iow6 = (~(Jcaiu6 | D7fpw6[12]));
assign Zeohu6 = (~(Q5iow6 & X5iow6));
assign X5iow6 = (~(Umhow6 & HRDATA[22]));
assign Q5iow6 = (~(Hrfpw6[6] & Qqhiu6));
assign Seohu6 = (~(E6iow6 & L6iow6));
assign L6iow6 = (~(Umhow6 & HRDATA[21]));
assign E6iow6 = (~(Hrfpw6[5] & Qqhiu6));
assign Leohu6 = (S6iow6 | Z6iow6);
assign Z6iow6 = (~(G7iow6 | Dk7ow6));
assign Dk7ow6 = (N7iow6 & S3kiu6);
assign S3kiu6 = (U7iow6 & B8iow6);
assign B8iow6 = (~(Toaiu6 & It2ju6));
assign U7iow6 = (Oe8ow6 | Cyfpw6[6]);
assign N7iow6 = (I8iow6 & Et0ju6);
assign I8iow6 = (~(L45iu6 & Llaow6));
assign S6iow6 = (Rk7ow6 ? S8fpw6[6] : P8iow6);
assign Rk7ow6 = (~(HREADY & W8iow6));
assign W8iow6 = (~(D9iow6 & K9iow6));
assign K9iow6 = (R9iow6 & Y9iow6);
assign Y9iow6 = (Faiow6 & Maiow6);
assign Maiow6 = (~(Taiow6 & N2ghu6));
assign Taiow6 = (~(D9oiu6 | Kq0iu6));
assign D9oiu6 = (!Whfiu6);
assign Faiow6 = (~(Abiow6 & Ae0iu6));
assign Abiow6 = (Pthiu6 & Mr0iu6);
assign R9iow6 = (Hbiow6 & Obiow6);
assign Obiow6 = (~(Vbiow6 & Xzmiu6));
assign Hbiow6 = (~(Hviiu6 & Gaziu6));
assign D9iow6 = (Cciow6 & T1jiu6);
assign T1jiu6 = (Jciow6 & Qciow6);
assign Qciow6 = (~(Us2ju6 & Yljiu6));
assign Jciow6 = (Xciow6 & Ediow6);
assign Ediow6 = (~(Ldiow6 & S6aiu6));
assign Ldiow6 = (~(Cyfpw6[0] | Cyfpw6[3]));
assign Xciow6 = (~(Zzniu6 & Qu7ow6));
assign Zzniu6 = (~(R2aiu6 | Mjfiu6));
assign Cciow6 = (Epjiu6 & Sdiow6);
assign Sdiow6 = (Wmaiu6 | Nloiu6);
assign Epjiu6 = (Zdiow6 & Geiow6);
assign Geiow6 = (Neiow6 & Ueiow6);
assign Ueiow6 = (Bfiow6 & Ifiow6);
assign Ifiow6 = (~(Lzhow6 & Raaow6));
assign Raaow6 = (Uyiiu6 & Uriiu6);
assign Lzhow6 = (Nbkiu6 & X1ziu6);
assign Bfiow6 = (E2ziu6 & Oe8ow6);
assign E2ziu6 = (~(Pfiow6 & Jjhiu6));
assign Neiow6 = (Wfiow6 & Dgiow6);
assign Dgiow6 = (~(Vviiu6 & Kgiow6));
assign Kgiow6 = (~(X1ziu6 & Rgiow6));
assign Rgiow6 = (D7fpw6[8] | D7fpw6[9]);
assign Vviiu6 = (Uyiiu6 & J9kiu6);
assign Wfiow6 = (~(Hviiu6 & Db0ju6));
assign Db0ju6 = (D7fpw6[10] & Tniiu6);
assign Hviiu6 = (Ygiow6 & J9kiu6);
assign Ygiow6 = (~(Lraiu6 | D7fpw6[14]));
assign Zdiow6 = (Fhiow6 & Mhiow6);
assign Mhiow6 = (Thiow6 & Aiiow6);
assign Aiiow6 = (~(Y31ju6 & Hiiow6));
assign Hiiow6 = (~(Oiiow6 & Viiow6));
assign Viiow6 = (N38ow6 | D7fpw6[15]);
assign Oiiow6 = (~(Cjiow6 | J1ziu6));
assign Cjiow6 = (Jjiow6 & P0piu6);
assign Jjiow6 = (~(Qjiow6 | O95iu6));
assign Thiow6 = (O4aiu6 | D7fpw6[3]);
assign Fhiow6 = (D0jiu6 & Veziu6);
assign Veziu6 = (B1aiu6 & Xjiow6);
assign Xjiow6 = (~(Y0jiu6 & Tfjiu6));
assign B1aiu6 = (!Ezhow6);
assign Ezhow6 = (O4oiu6 & Taaiu6);
assign D0jiu6 = (Ekiow6 & Lkiow6);
assign Lkiow6 = (Skiow6 & Zkiow6);
assign Zkiow6 = (~(Gliow6 & Nliow6));
assign Nliow6 = (~(Qxoiu6 | D7fpw6[13]));
assign Gliow6 = (J9kiu6 & Q5aiu6);
assign Skiow6 = (~(De6ow6 & F9aju6));
assign Ekiow6 = (Uliow6 & Bmiow6);
assign Bmiow6 = (~(Evyiu6 & W0piu6));
assign W0piu6 = (~(Ftjiu6 | Lraiu6));
assign Evyiu6 = (Mtjiu6 & X1ziu6);
assign Uliow6 = (O4aiu6 | Cyfpw6[0]);
assign O4aiu6 = (~(Nu9ow6 & K9aiu6));
assign Nu9ow6 = (Imiow6 & Pmiow6);
assign Pmiow6 = (~(D7fpw6[14] | Cyfpw6[3]));
assign Imiow6 = (Ya1ju6 & Hzziu6);
assign P8iow6 = (~(Wmiow6 & Dniow6));
assign Dniow6 = (Ad8iu6 | Hm7ow6);
assign Hm7ow6 = (~(Zlhow6 | Th2ju6));
assign Zlhow6 = (~(Kniow6 & Rniow6));
assign Rniow6 = (Yniow6 & Foiow6);
assign Foiow6 = (Hujiu6 | I6jiu6);
assign Yniow6 = (Moiow6 & S4jiu6);
assign S4jiu6 = (~(Toiow6 & Ia8iu6));
assign Toiow6 = (~(C27ow6 | Ftjiu6));
assign C27ow6 = (!Wliiu6);
assign Moiow6 = (~(J1ziu6 & Ia8iu6));
assign J1ziu6 = (Wliiu6 & D7fpw6[11]);
assign Wliiu6 = (Mtjiu6 & Gaziu6);
assign Gaziu6 = (!D7fpw6[13]);
assign Kniow6 = (Ubkiu6 & Apiow6);
assign Apiow6 = (E4jiu6 | Ae0iu6);
assign Ubkiu6 = (Ymiiu6 & Hpiow6);
assign Hpiow6 = (Hujiu6 | Aujiu6);
assign Hujiu6 = (!Th2ju6);
assign Th2ju6 = (Xiiiu6 & Kxziu6);
assign Ymiiu6 = (Xl0ju6 | Qpaju6);
assign Qpaju6 = (!Kxziu6);
assign Xl0ju6 = (!R7jiu6);
assign Wmiow6 = (Dzjiu6 | Cn7ow6);
assign Cn7ow6 = (Opiow6 & Oaiiu6);
assign Oaiiu6 = (~(Vpiow6 & J9kiu6));
assign Vpiow6 = (~(Co6ow6 | Ae0iu6));
assign Opiow6 = (~(Ia8iu6 & Ozziu6));
assign Eeohu6 = (~(Cqiow6 & Jqiow6));
assign Jqiow6 = (~(Umhow6 & HRDATA[20]));
assign Cqiow6 = (~(Hrfpw6[4] & Qqhiu6));
assign Xdohu6 = (Eh6iu6 ? Sufpw6[0] : Qqiow6);
assign Qqiow6 = (Xqiow6 & Ophiu6);
assign Xqiow6 = (N6piu6 | Sufpw6[1]);
assign Qdohu6 = (Eh6iu6 ? L3ehu6 : Fnpiu6);
assign Fnpiu6 = (!Ejpiu6);
assign Jdohu6 = (~(Eriow6 & Lriow6));
assign Lriow6 = (Sriow6 & Zriow6);
assign Zriow6 = (~(Egziu6 & Eafpw6[11]));
assign Sriow6 = (Gsiow6 & Sgziu6);
assign Gsiow6 = (~(Zgziu6 & Uumiu6));
assign Uumiu6 = (~(Nsiow6 & Usiow6));
assign Usiow6 = (Btiow6 & Itiow6);
assign Itiow6 = (Tgcow6 | Pkdow6);
assign Tgcow6 = (Ptiow6 & Wtiow6);
assign Wtiow6 = (Duiow6 & Kuiow6);
assign Kuiow6 = (~(Dyeow6 & Re4ju6));
assign Duiow6 = (Iydow6 | Uosiu6);
assign Uosiu6 = (Ruiow6 & Yuiow6);
assign Yuiow6 = (Fviow6 & Mviow6);
assign Mviow6 = (~(Tzfpw6[11] & Yvgiu6));
assign Fviow6 = (Tviow6 & Awiow6);
assign Awiow6 = (~(F0eow6 & Vbgpw6[11]));
assign Tviow6 = (~(Odgpw6[11] & M0eow6));
assign Ruiow6 = (Hwiow6 & Owiow6);
assign Owiow6 = (~(Bagpw6[11] & M6eiu6));
assign Hwiow6 = (~(STCALIB[11] & H1eow6));
assign Ptiow6 = (Vwiow6 & Cxiow6);
assign Cxiow6 = (~(Qtfow6 & Ag4ju6));
assign Vwiow6 = (~(HRDATA[11] & Q2eow6));
assign Btiow6 = (Jxiow6 & Dldow6);
assign Jxiow6 = (Kfcow6 | Uqdow6);
assign Kfcow6 = (Qxiow6 & Xxiow6);
assign Xxiow6 = (Eyiow6 & Lyiow6);
assign Lyiow6 = (~(Dyeow6 & Jw3ju6));
assign Eyiow6 = (Iydow6 | Tmqiu6);
assign Tmqiu6 = (Syiow6 & Zyiow6);
assign Zyiow6 = (Gziow6 & Nziow6);
assign Nziow6 = (Uziow6 & B0jow6);
assign Uziow6 = (~(STCALIB[3] & H1eow6));
assign Gziow6 = (I0jow6 & P0jow6);
assign P0jow6 = (~(Odgpw6[3] & M0eow6));
assign I0jow6 = (~(Tzfpw6[3] & Yvgiu6));
assign Syiow6 = (W0jow6 & D1jow6);
assign D1jow6 = (K1jow6 & R1jow6);
assign R1jow6 = (~(Bagpw6[3] & M6eiu6));
assign K1jow6 = (~(F0eow6 & Vbgpw6[3]));
assign W0jow6 = (Y1jow6 & F2jow6);
assign F2jow6 = (Qkgiu6 | Ngfiu6);
assign Y1jow6 = (~(ECOREVNUM[3] & I5eow6));
assign Qxiow6 = (M2jow6 & T2jow6);
assign T2jow6 = (~(Qtfow6 & Lx3ju6));
assign M2jow6 = (~(HRDATA[3] & Q2eow6));
assign Nsiow6 = (A3jow6 & H3jow6);
assign H3jow6 = (Ahcow6 | Kldow6);
assign Ahcow6 = (O3jow6 & V3jow6);
assign V3jow6 = (C4jow6 & J4jow6);
assign J4jow6 = (Rcfow6 | C34ju6);
assign C4jow6 = (Iydow6 | U8uiu6);
assign U8uiu6 = (Q4jow6 & X4jow6);
assign X4jow6 = (E5jow6 & L5jow6);
assign L5jow6 = (~(STCALIB[19] & H1eow6));
assign E5jow6 = (S5jow6 & Z5jow6);
assign Z5jow6 = (~(Tzfpw6[19] & Yvgiu6));
assign S5jow6 = (~(Bagpw6[19] & M6eiu6));
assign Q4jow6 = (~(G6jow6 | I5eow6));
assign G6jow6 = (~(N6jow6 & U6jow6));
assign U6jow6 = (~(Odgpw6[19] & M0eow6));
assign N6jow6 = (~(F0eow6 & Vbgpw6[19]));
assign O3jow6 = (B7jow6 & I7jow6);
assign I7jow6 = (~(Qtfow6 & L44ju6));
assign B7jow6 = (~(HRDATA[19] & Q2eow6));
assign A3jow6 = (Yfcow6 | Spdow6);
assign Yfcow6 = (P7jow6 & W7jow6);
assign W7jow6 = (Iydow6 | Wtviu6);
assign Wtviu6 = (D8jow6 & K8jow6);
assign K8jow6 = (~(F0eow6 & Vbgpw6[27]));
assign D8jow6 = (R8jow6 & Yreow6);
assign R8jow6 = (~(Odgpw6[27] & M0eow6));
assign P7jow6 = (Y8jow6 & F9jow6);
assign F9jow6 = (~(C2eow6 & M9jow6));
assign M9jow6 = (~(O94ju6 & T9jow6));
assign T9jow6 = (Aajow6 | Bz3ju6);
assign O94ju6 = (~(Hajow6 & Oajow6));
assign Oajow6 = (Vajow6 | J2eow6);
assign Hajow6 = (Cbjow6 & Aajow6);
assign Aajow6 = (~(Jbjow6 & Qbjow6));
assign Cbjow6 = (~(Xbjow6 & Ecjow6));
assign Xbjow6 = (J2eow6 & Lcjow6);
assign Y8jow6 = (~(HRDATA[27] & Q2eow6));
assign Eriow6 = (Scjow6 & Zcjow6);
assign Zcjow6 = (~(Zsfpw6[10] & Cmziu6));
assign Scjow6 = (~(vis_pc_o[10] & Jmziu6));
assign Cdohu6 = (~(Gdjow6 & Ndjow6));
assign Ndjow6 = (Udjow6 & Bejow6);
assign Bejow6 = (~(Egziu6 & Eafpw6[9]));
assign Udjow6 = (Iejow6 & Sgziu6);
assign Iejow6 = (~(Zgziu6 & S0niu6));
assign S0niu6 = (~(Pejow6 & Wejow6));
assign Wejow6 = (Dfjow6 & Kfjow6);
assign Kfjow6 = (~(Mmdow6 & Ew6ow6));
assign Ew6ow6 = (~(Rfjow6 & Yfjow6));
assign Yfjow6 = (Fgjow6 & Mgjow6);
assign Mgjow6 = (Rcfow6 | Mu3ju6);
assign Mu3ju6 = (Tgjow6 & Ahjow6);
assign Ahjow6 = (Hhjow6 & Ohjow6);
assign Ohjow6 = (Rqfow6 | I40iu6);
assign Hhjow6 = (Ipfow6 | B40iu6);
assign Tgjow6 = (Vhjow6 & Cijow6);
assign Cijow6 = (Ppfow6 | W40iu6);
assign Vhjow6 = (Kqfow6 | P40iu6);
assign Fgjow6 = (Iydow6 | Ovpiu6);
assign Ovpiu6 = (Jijow6 & Qijow6);
assign Qijow6 = (Xijow6 & Ejjow6);
assign Ejjow6 = (Ljjow6 & Sjjow6);
assign Sjjow6 = (~(Odgpw6[1] & M0eow6));
assign Ljjow6 = (Zjjow6 & Gkjow6);
assign Gkjow6 = (~(Fpgiu6 & Qqdhu6));
assign Zjjow6 = (~(Tzfpw6[1] & Yvgiu6));
assign Xijow6 = (Nkjow6 & Ukjow6);
assign Ukjow6 = (~(ECOREVNUM[1] & I5eow6));
assign Nkjow6 = (~(Y5eiu6 & Dvghu6));
assign Jijow6 = (Bljow6 & Iljow6);
assign Iljow6 = (Pljow6 & Wljow6);
assign Wljow6 = (~(F0eow6 & Vbgpw6[1]));
assign Pljow6 = (~(Bagpw6[1] & M6eiu6));
assign Bljow6 = (Dmjow6 & Kmjow6);
assign Kmjow6 = (~(STCALIB[1] & H1eow6));
assign Dmjow6 = (Qkgiu6 | Siciu6);
assign Rfjow6 = (Rmjow6 & Ymjow6);
assign Ymjow6 = (~(Qtfow6 & Ex3ju6));
assign Ex3ju6 = (~(Fnjow6 & Mnjow6));
assign Mnjow6 = (Tnjow6 & Aojow6);
assign Aojow6 = (Kqfow6 | F60iu6);
assign Tnjow6 = (Ipfow6 | D50iu6);
assign Fnjow6 = (Hojow6 & Oojow6);
assign Oojow6 = (Rqfow6 | K50iu6);
assign Hojow6 = (Ppfow6 | E90iu6);
assign Rmjow6 = (~(HRDATA[1] & Q2eow6));
assign Dfjow6 = (Vojow6 & Dldow6);
assign Vojow6 = (Pkdow6 | Xv6ow6);
assign Xv6ow6 = (Cpjow6 & Jpjow6);
assign Jpjow6 = (Qpjow6 & Xpjow6);
assign Xpjow6 = (Rcfow6 | Uc4ju6);
assign Uc4ju6 = (Eqjow6 & Lqjow6);
assign Lqjow6 = (Sqjow6 & Zqjow6);
assign Zqjow6 = (Ipfow6 | Ga0iu6);
assign Sqjow6 = (Ppfow6 | Bb0iu6);
assign Eqjow6 = (Grjow6 & Nrjow6);
assign Nrjow6 = (Kqfow6 | Ua0iu6);
assign Grjow6 = (Rqfow6 | Na0iu6);
assign Qpjow6 = (Iydow6 | Ibsiu6);
assign Ibsiu6 = (Urjow6 & Bsjow6);
assign Bsjow6 = (Isjow6 & Psjow6);
assign Psjow6 = (Wsjow6 & B0jow6);
assign B0jow6 = (~(Rzciu6 & Dtjow6));
assign Wsjow6 = (~(Bagpw6[9] & M6eiu6));
assign Isjow6 = (Ktjow6 & Rtjow6);
assign Rtjow6 = (~(Tzfpw6[9] & Yvgiu6));
assign Ktjow6 = (~(F0eow6 & Vbgpw6[9]));
assign Urjow6 = (Ytjow6 & Qgeow6);
assign Ytjow6 = (Fujow6 & Mujow6);
assign Mujow6 = (~(STCALIB[9] & H1eow6));
assign Fujow6 = (~(M0eow6 & Odgpw6[9]));
assign Cpjow6 = (Tujow6 & Avjow6);
assign Avjow6 = (~(Qtfow6 & Hg4ju6));
assign Hg4ju6 = (~(Hvjow6 & Ovjow6));
assign Ovjow6 = (Vvjow6 & Cwjow6);
assign Cwjow6 = (Rqfow6 | Pb0iu6);
assign Vvjow6 = (Ppfow6 | U30iu6);
assign Hvjow6 = (Jwjow6 & Qwjow6);
assign Qwjow6 = (Kqfow6 | Wb0iu6);
assign Jwjow6 = (Ipfow6 | Ib0iu6);
assign Tujow6 = (~(HRDATA[9] & Q2eow6));
assign Pejow6 = (Xwjow6 & Exjow6);
assign Exjow6 = (~(Fmdow6 & Cv6ow6));
assign Cv6ow6 = (~(Lxjow6 & Sxjow6));
assign Sxjow6 = (Iydow6 | Wfviu6);
assign Wfviu6 = (Zxjow6 & Gyjow6);
assign Gyjow6 = (~(F0eow6 & Vbgpw6[25]));
assign Zxjow6 = (Nyjow6 & Yreow6);
assign Nyjow6 = (~(M0eow6 & Odgpw6[25]));
assign Lxjow6 = (Uyjow6 & Bzjow6);
assign Bzjow6 = (~(C2eow6 & Izjow6));
assign Izjow6 = (~(Pzjow6 & Wzjow6));
assign Wzjow6 = (D0kow6 | Bz3ju6);
assign Pzjow6 = (~(M84ju6 & K0kow6));
assign K0kow6 = (V94ju6 | Hv3ju6);
assign V94ju6 = (~(R0kow6 & Y0kow6));
assign Y0kow6 = (F1kow6 & M1kow6);
assign M1kow6 = (Ipfow6 | T60iu6);
assign F1kow6 = (Ppfow6 | O70iu6);
assign R0kow6 = (T1kow6 & A2kow6);
assign A2kow6 = (Kqfow6 | H70iu6);
assign T1kow6 = (Rqfow6 | A70iu6);
assign M84ju6 = (H2kow6 & D0kow6);
assign D0kow6 = (~(O2kow6 & Jbjow6));
assign O2kow6 = (Sveow6 ? V2kow6 : Qbjow6);
assign Sveow6 = (C3kow6 | Gweow6);
assign H2kow6 = (~(Nweow6 & Hv3ju6));
assign Nweow6 = (J3kow6 & Q3kow6);
assign Q3kow6 = (X3kow6 & E4kow6);
assign E4kow6 = (Ipfow6 | Dc0iu6);
assign X3kow6 = (Rqfow6 | R50iu6);
assign J3kow6 = (L4kow6 & S4kow6);
assign S4kow6 = (Ppfow6 | M60iu6);
assign L4kow6 = (Kqfow6 | Y50iu6);
assign Uyjow6 = (~(HRDATA[25] & Q2eow6));
assign Xwjow6 = (Kldow6 | Ou6ow6);
assign Ou6ow6 = (Z4kow6 & G5kow6);
assign G5kow6 = (N5kow6 & U5kow6);
assign U5kow6 = (Rcfow6 | F14ju6);
assign F14ju6 = (B6kow6 & I6kow6);
assign I6kow6 = (P6kow6 & W6kow6);
assign W6kow6 = (Ipfow6 | V70iu6);
assign P6kow6 = (Rqfow6 | C80iu6);
assign B6kow6 = (D7kow6 & K7kow6);
assign K7kow6 = (Ppfow6 | Q80iu6);
assign D7kow6 = (Kqfow6 | J80iu6);
assign N5kow6 = (Iydow6 | Nutiu6);
assign Nutiu6 = (R7kow6 & Y7kow6);
assign Y7kow6 = (F8kow6 & M8kow6);
assign M8kow6 = (~(Tzfpw6[17] & Yvgiu6));
assign F8kow6 = (T8kow6 & A9kow6);
assign A9kow6 = (W6ciu6 | Qkgiu6);
assign W6ciu6 = (~(H9kow6 & Ydeow6));
assign H9kow6 = (~(Feeow6 | E2fow6));
assign T8kow6 = (~(Odgpw6[17] & M0eow6));
assign R7kow6 = (O9kow6 & V9kow6);
assign V9kow6 = (~(F0eow6 & Vbgpw6[17]));
assign O9kow6 = (Cakow6 & Jakow6);
assign Jakow6 = (~(STCALIB[17] & H1eow6));
assign Cakow6 = (~(Bagpw6[17] & M6eiu6));
assign Z4kow6 = (Qakow6 & Xakow6);
assign Xakow6 = (~(Qtfow6 & Ff4ju6));
assign Ff4ju6 = (~(Ebkow6 & Lbkow6));
assign Lbkow6 = (Sbkow6 & Zbkow6);
assign Zbkow6 = (Ipfow6 | X80iu6);
assign Sbkow6 = (Rqfow6 | L90iu6);
assign Ebkow6 = (Gckow6 & Nckow6);
assign Nckow6 = (Ppfow6 | Z90iu6);
assign Gckow6 = (Kqfow6 | S90iu6);
assign Qakow6 = (~(HRDATA[17] & Q2eow6));
assign Gdjow6 = (Uckow6 & Bdkow6);
assign Bdkow6 = (~(Zsfpw6[8] & Cmziu6));
assign Uckow6 = (~(vis_pc_o[8] & Jmziu6));
assign Vcohu6 = (~(Idkow6 & Pdkow6));
assign Pdkow6 = (Wdkow6 & Dekow6);
assign Dekow6 = (~(Egziu6 & Eafpw6[15]));
assign Wdkow6 = (Kekow6 & Sgziu6);
assign Kekow6 = (Ft6ow6 | Ggmiu6);
assign Ggmiu6 = (Rekow6 & Yekow6);
assign Yekow6 = (Ffkow6 & Mfkow6);
assign Mfkow6 = (H78ow6 | Kldow6);
assign Ffkow6 = (Tfkow6 & Dldow6);
assign Tfkow6 = (~(Mmdow6 & X88ow6));
assign Rekow6 = (Agkow6 & Hgkow6);
assign Hgkow6 = (~(V78ow6 & Fmdow6));
assign Agkow6 = (Q88ow6 | Pkdow6);
assign Idkow6 = (Ogkow6 & Vgkow6);
assign Vgkow6 = (~(Zsfpw6[14] & Cmziu6));
assign Ogkow6 = (~(vis_pc_o[14] & Jmziu6));
assign Ocohu6 = (~(Chkow6 & Jhkow6));
assign Jhkow6 = (Qhkow6 & Xhkow6);
assign Xhkow6 = (~(Zsfpw6[21] & Cmziu6));
assign Qhkow6 = (Eikow6 & Likow6);
assign Likow6 = (Ft6ow6 | Nvliu6);
assign Nvliu6 = (Sikow6 & Zikow6);
assign Zikow6 = (Gjkow6 & Njkow6);
assign Njkow6 = (G6cow6 | Eccow6);
assign G6cow6 = (Ujkow6 & Bkkow6);
assign Bkkow6 = (Ikkow6 & Pkkow6);
assign Pkkow6 = (Rcfow6 | Wkkow6);
assign Wkkow6 = (!O24ju6);
assign Ikkow6 = (Iydow6 | Ntuiu6);
assign Ntuiu6 = (Dlkow6 & Klkow6);
assign Klkow6 = (Rlkow6 & Ylkow6);
assign Ylkow6 = (Fmkow6 & Mmkow6);
assign Mmkow6 = (Tmkow6 & Ankow6);
assign Ankow6 = (~(Odgpw6[22] & M0eow6));
assign Tmkow6 = (~(STCALIB[22] & H1eow6));
assign Fmkow6 = (Hnkow6 & Onkow6);
assign Onkow6 = (~(Tzdiu6 & R4gpw6[4]));
assign Hnkow6 = (~(I3fiu6 & R4gpw6[12]));
assign Rlkow6 = (Vnkow6 & Cokow6);
assign Cokow6 = (Jokow6 & Qokow6);
assign Qokow6 = (~(Tzfpw6[22] & Yvgiu6));
assign Jokow6 = (~(Hqgiu6 & L1gpw6[0]));
assign Vnkow6 = (Xokow6 & Epkow6);
assign Epkow6 = (~(S1fiu6 & R4gpw6[36]));
assign Xokow6 = (~(G2fiu6 & R4gpw6[28]));
assign Dlkow6 = (Lpkow6 & Spkow6);
assign Spkow6 = (Zpkow6 & Gqkow6);
assign Gqkow6 = (Nqkow6 & Uqkow6);
assign Uqkow6 = (~(C0fiu6 & R4gpw6[60]));
assign Nqkow6 = (~(F0eow6 & Vbgpw6[22]));
assign Zpkow6 = (Brkow6 & Irkow6);
assign Irkow6 = (~(Bagpw6[22] & M6eiu6));
assign Brkow6 = (~(E1fiu6 & R4gpw6[44]));
assign Lpkow6 = (Prkow6 & Wrkow6);
assign Wrkow6 = (~(T7eow6 & Dskow6));
assign Dskow6 = (~(Kskow6 & Rskow6));
assign Rskow6 = (Yskow6 & Ftkow6);
assign Ftkow6 = (Mtkow6 & Ttkow6);
assign Ttkow6 = (Aukow6 & Hukow6);
assign Hukow6 = (~(Odgpw6[8] | Odgpw6[9]));
assign Aukow6 = (~(Odgpw6[6] | Odgpw6[7]));
assign Mtkow6 = (Oukow6 & Vukow6);
assign Vukow6 = (~(Odgpw6[4] | Odgpw6[5]));
assign Oukow6 = (~(Odgpw6[31] | Odgpw6[3]));
assign Yskow6 = (Cvkow6 & Jvkow6);
assign Jvkow6 = (Qvkow6 & Xvkow6);
assign Xvkow6 = (~(Odgpw6[2] | Odgpw6[30]));
assign Qvkow6 = (~(Odgpw6[28] | Odgpw6[29]));
assign Cvkow6 = (Ewkow6 & Lwkow6);
assign Lwkow6 = (~(Odgpw6[26] | Odgpw6[27]));
assign Ewkow6 = (~(Odgpw6[24] | Odgpw6[25]));
assign Kskow6 = (Swkow6 & Zwkow6);
assign Zwkow6 = (Gxkow6 & Nxkow6);
assign Nxkow6 = (Uxkow6 & Bykow6);
assign Bykow6 = (~(Odgpw6[22] | Odgpw6[23]));
assign Uxkow6 = (~(Odgpw6[20] | Odgpw6[21]));
assign Gxkow6 = (Iykow6 & Pykow6);
assign Pykow6 = (~(Odgpw6[19] | Odgpw6[1]));
assign Iykow6 = (~(Odgpw6[17] | Odgpw6[18]));
assign Swkow6 = (Wykow6 & Dzkow6);
assign Dzkow6 = (Kzkow6 & Rzkow6);
assign Rzkow6 = (~(Odgpw6[15] | Odgpw6[16]));
assign Kzkow6 = (~(Odgpw6[13] | Odgpw6[14]));
assign Wykow6 = (Yzkow6 & F0low6);
assign F0low6 = (~(Odgpw6[11] | Odgpw6[12]));
assign Yzkow6 = (~(Odgpw6[0] | Odgpw6[10]));
assign Prkow6 = (M0low6 & T0low6);
assign T0low6 = (~(Q0fiu6 & R4gpw6[52]));
assign M0low6 = (~(U2fiu6 & R4gpw6[20]));
assign Ujkow6 = (A1low6 & H1low6);
assign H1low6 = (Uafow6 | R04ju6);
assign A1low6 = (~(HRDATA[22] & Q2eow6));
assign Gjkow6 = (L5cow6 | Vacow6);
assign Vacow6 = (O1low6 & Dtcow6);
assign L5cow6 = (V1low6 & C2low6);
assign C2low6 = (J2low6 & Q2low6);
assign Q2low6 = (~(Dyeow6 & Ye4ju6));
assign J2low6 = (Iydow6 | N9tiu6);
assign N9tiu6 = (X2low6 & E3low6);
assign E3low6 = (L3low6 & S3low6);
assign S3low6 = (Z3low6 & G4low6);
assign G4low6 = (N4low6 & U4low6);
assign U4low6 = (~(Tzdiu6 & R4gpw6[2]));
assign N4low6 = (~(S1fiu6 & R4gpw6[34]));
assign Z3low6 = (B5low6 & I5low6);
assign I5low6 = (~(STCALIB[14] & H1eow6));
assign B5low6 = (~(F0eow6 & Vbgpw6[14]));
assign L3low6 = (P5low6 & W5low6);
assign W5low6 = (D6low6 & K6low6);
assign K6low6 = (~(U2fiu6 & R4gpw6[18]));
assign D6low6 = (~(I3fiu6 & R4gpw6[10]));
assign P5low6 = (R6low6 & Y6low6);
assign Y6low6 = (U5ciu6 | Qkgiu6);
assign U5ciu6 = (~(Ydeow6 & F7low6));
assign F7low6 = (~(Okgow6 & M7low6));
assign M7low6 = (~(T7low6 & A8low6));
assign T7low6 = (~(H8low6 & O8low6));
assign H8low6 = (E2fow6 ? C9low6 : V8low6);
assign C9low6 = (~(Z2fow6 | J9low6));
assign J9low6 = (~(B4fow6 | Nggow6));
assign V8low6 = (F6fow6 & Q9low6);
assign Q9low6 = (H7fow6 | Hdgow6);
assign R6low6 = (~(Q0fiu6 & R4gpw6[50]));
assign X2low6 = (X9low6 & Ealow6);
assign Ealow6 = (Lalow6 & Salow6);
assign Salow6 = (Zalow6 & Gblow6);
assign Gblow6 = (~(Tzfpw6[14] & Yvgiu6));
assign Zalow6 = (~(Odgpw6[14] & M0eow6));
assign Lalow6 = (Nblow6 & Ublow6);
assign Ublow6 = (~(C0fiu6 & R4gpw6[58]));
assign Nblow6 = (~(E1fiu6 & R4gpw6[42]));
assign X9low6 = (Bclow6 & Qgeow6);
assign Bclow6 = (Iclow6 & Pclow6);
assign Pclow6 = (~(Bagpw6[14] & M6eiu6));
assign Iclow6 = (~(G2fiu6 & R4gpw6[26]));
assign V1low6 = (Wclow6 & Ddlow6);
assign Ddlow6 = (Uafow6 | Id4ju6);
assign Wclow6 = (~(HRDATA[14] & Q2eow6));
assign Sikow6 = (Kdlow6 & Rdlow6);
assign Rdlow6 = (~(X4cow6 & Cbcow6));
assign Cbcow6 = (~(Ydlow6 & W9how6));
assign X4cow6 = (~(Felow6 & Melow6));
assign Melow6 = (Iydow6 | Bewiu6);
assign Bewiu6 = (Telow6 & Aflow6);
assign Aflow6 = (Hflow6 & Oflow6);
assign Oflow6 = (Vflow6 & Cglow6);
assign Cglow6 = (Jglow6 & Qglow6);
assign Qglow6 = (~(Odgpw6[30] & M0eow6));
assign Jglow6 = (Tpgiu6 | Xglow6);
assign Vflow6 = (Ehlow6 & Lhlow6);
assign Lhlow6 = (~(E1fiu6 & R4gpw6[46]));
assign Ehlow6 = (~(Tzdiu6 & R4gpw6[6]));
assign Hflow6 = (Shlow6 & Zhlow6);
assign Zhlow6 = (~(U2fiu6 & R4gpw6[22]));
assign Shlow6 = (Gilow6 & Nilow6);
assign Nilow6 = (~(STCALIB[24] & H1eow6));
assign Gilow6 = (~(G2fiu6 & R4gpw6[30]));
assign Telow6 = (Uilow6 & Bjlow6);
assign Bjlow6 = (Ijlow6 & Pjlow6);
assign Pjlow6 = (Wjlow6 & Dklow6);
assign Dklow6 = (~(Hqgiu6 & H8gpw6[0]));
assign Wjlow6 = (~(I3fiu6 & R4gpw6[14]));
assign Ijlow6 = (Kklow6 & Rklow6);
assign Rklow6 = (~(C0fiu6 & R4gpw6[62]));
assign Kklow6 = (~(S1fiu6 & R4gpw6[38]));
assign Uilow6 = (Yklow6 & Qgeow6);
assign Yklow6 = (Fllow6 & Mllow6);
assign Mllow6 = (~(Q0fiu6 & R4gpw6[54]));
assign Fllow6 = (~(Pceow6 & Tllow6));
assign Tllow6 = (Nzhiu6 | Vbgpw6[30]);
assign Felow6 = (Amlow6 & Hmlow6);
assign Hmlow6 = (~(C2eow6 & Omlow6));
assign Omlow6 = (~(Vmlow6 & A94ju6));
assign A94ju6 = (~(Cnlow6 & Jnlow6));
assign Jnlow6 = (~(Qnlow6 & Queow6));
assign Qnlow6 = (Xnlow6 & Zveow6);
assign Xnlow6 = (Azfow6 | Kqfow6);
assign Cnlow6 = (J2eow6 ? Eolow6 : Zx3ju6);
assign Vmlow6 = (~(Lolow6 & Vh3ju6));
assign Lolow6 = (Queow6 & Zveow6);
assign Zveow6 = (Solow6 | C3kow6);
assign Amlow6 = (~(HRDATA[30] & Q2eow6));
assign Kdlow6 = (~(Xbcow6 & N6cow6));
assign N6cow6 = (~(Zolow6 & Gplow6));
assign Gplow6 = (Nplow6 & Uplow6);
assign Uplow6 = (~(Dyeow6 & Og4ju6));
assign Nplow6 = (Iydow6 | Kkriu6);
assign Kkriu6 = (Bqlow6 & Iqlow6);
assign Iqlow6 = (Pqlow6 & Wqlow6);
assign Wqlow6 = (Drlow6 & Krlow6);
assign Krlow6 = (Rrlow6 & Yrlow6);
assign Yrlow6 = (~(Odgpw6[6] & M0eow6));
assign Rrlow6 = (~(Q0fiu6 & R4gpw6[48]));
assign Drlow6 = (Fslow6 & Mslow6);
assign Mslow6 = (~(Bagpw6[6] & M6eiu6));
assign Fslow6 = (~(C0fiu6 & R4gpw6[56]));
assign Pqlow6 = (Tslow6 & Atlow6);
assign Atlow6 = (~(E1fiu6 & R4gpw6[40]));
assign Tslow6 = (Htlow6 & Otlow6);
assign Otlow6 = (~(Tzfpw6[6] & Yvgiu6));
assign Htlow6 = (~(STCALIB[6] & H1eow6));
assign Bqlow6 = (Vtlow6 & Culow6);
assign Culow6 = (Julow6 & Qulow6);
assign Qulow6 = (~(F0eow6 & Vbgpw6[6]));
assign Julow6 = (Xulow6 & Evlow6);
assign Evlow6 = (~(S1fiu6 & R4gpw6[32]));
assign Xulow6 = (~(G2fiu6 & R4gpw6[24]));
assign Vtlow6 = (Lvlow6 & Svlow6);
assign Svlow6 = (~(U2fiu6 & R4gpw6[16]));
assign Lvlow6 = (Zvlow6 & Gwlow6);
assign Gwlow6 = (~(I3fiu6 & R4gpw6[8]));
assign Zvlow6 = (~(Tzdiu6 & R4gpw6[0]));
assign Zolow6 = (Nwlow6 & Uwlow6);
assign Uwlow6 = (Uafow6 | Yt3ju6);
assign Uafow6 = (!Qtfow6);
assign Nwlow6 = (~(HRDATA[6] & Q2eow6));
assign Xbcow6 = (~(K3how6 | Df3ju6));
assign Eikow6 = (~(Egziu6 & Eafpw6[22]));
assign Chkow6 = (Lccow6 & Bxlow6);
assign Bxlow6 = (~(vis_pc_o[21] & Jmziu6));
assign Lccow6 = (Sgziu6 & Ixlow6);
assign Ixlow6 = (Svkiu6 | Ft6ow6);
assign Ft6ow6 = (!Zgziu6);
assign Svkiu6 = (~(Pxlow6 & Ytcow6));
assign Ytcow6 = (Wxlow6 & H5how6);
assign Wxlow6 = (Tucow6 ? Oh3ju6 : Dylow6);
assign Oh3ju6 = (Kylow6 & Kf3ju6);
assign Kylow6 = (L7how6 | Df3ju6);
assign Dylow6 = (~(Rylow6 & Yylow6));
assign Yylow6 = (~(Fzlow6 & C0ehu6));
assign Fzlow6 = (Pthiu6 & Cyfpw6[5]);
assign Rylow6 = (C6how6 & Mzlow6);
assign Pxlow6 = (Ydlow6 & Tzlow6);
assign Ydlow6 = (Avcow6 | Ktcow6);
assign Hcohu6 = (~(A0mow6 & H0mow6));
assign H0mow6 = (O0mow6 & V0mow6);
assign V0mow6 = (~(Egziu6 & Eafpw6[10]));
assign Egziu6 = (Ar8iu6 & Et8iu6);
assign O0mow6 = (C1mow6 & Sgziu6);
assign Sgziu6 = (~(Ar8iu6 & J1mow6));
assign J1mow6 = (~(Q1mow6 & X1mow6));
assign X1mow6 = (~(Jydhu6 & Zmfiu6));
assign Zmfiu6 = (!Emfiu6);
assign Q1mow6 = (E2mow6 & Dp8iu6);
assign E2mow6 = (~(Qwdhu6 & M2biu6));
assign Ar8iu6 = (!Jmziu6);
assign C1mow6 = (~(Zgziu6 & Oymiu6));
assign Oymiu6 = (~(L2mow6 & S2mow6));
assign S2mow6 = (Z2mow6 & G3mow6);
assign G3mow6 = (Plcow6 | Pkdow6);
assign Pkdow6 = (Eccow6 & N3mow6);
assign N3mow6 = (~(Ktcow6 & U3mow6));
assign U3mow6 = (~(B4mow6 & I4mow6));
assign I4mow6 = (~(P4mow6 & Yahow6));
assign P4mow6 = (E6oiu6 | W4mow6);
assign W4mow6 = (F9aju6 & Nlaiu6);
assign E6oiu6 = (Cyfpw6[3] & Tr0iu6);
assign B4mow6 = (~(Jdhow6 | K2aiu6));
assign Jdhow6 = (T23ju6 & Cyfpw6[3]);
assign T23ju6 = (~(Tfjiu6 | Tr0iu6));
assign Eccow6 = (Tzlow6 & D5mow6);
assign D5mow6 = (!Ovcow6);
assign Ovcow6 = (Ktcow6 & K5mow6);
assign K5mow6 = (~(C0ehu6 & R5mow6));
assign R5mow6 = (~(G7oiu6 & Y5mow6));
assign Y5mow6 = (Y2oiu6 | Tr0iu6);
assign Plcow6 = (F6mow6 & M6mow6);
assign M6mow6 = (T6mow6 & A7mow6);
assign A7mow6 = (Rcfow6 | Id4ju6);
assign Id4ju6 = (H7mow6 & O7mow6);
assign O7mow6 = (V7mow6 & C8mow6);
assign C8mow6 = (Ipfow6 | Z90iu6);
assign V7mow6 = (Kqfow6 | Na0iu6);
assign H7mow6 = (J8mow6 & Q8mow6);
assign Q8mow6 = (Rqfow6 | Ga0iu6);
assign J8mow6 = (Ppfow6 | Ua0iu6);
assign T6mow6 = (Iydow6 | Bisiu6);
assign Bisiu6 = (X8mow6 & E9mow6);
assign E9mow6 = (L9mow6 & S9mow6);
assign S9mow6 = (~(Tzfpw6[10] & Yvgiu6));
assign L9mow6 = (Z9mow6 & Gamow6);
assign Gamow6 = (~(F0eow6 & Vbgpw6[10]));
assign Z9mow6 = (~(Odgpw6[10] & M0eow6));
assign X8mow6 = (Namow6 & Uamow6);
assign Uamow6 = (~(Bagpw6[10] & M6eiu6));
assign Namow6 = (~(STCALIB[10] & H1eow6));
assign F6mow6 = (Bbmow6 & Ibmow6);
assign Ibmow6 = (~(Qtfow6 & Og4ju6));
assign Og4ju6 = (~(Pbmow6 & Wbmow6));
assign Wbmow6 = (Dcmow6 & Kcmow6);
assign Kcmow6 = (Kqfow6 | Pb0iu6);
assign Dcmow6 = (Ppfow6 | Wb0iu6);
assign Pbmow6 = (Rcmow6 & Ycmow6);
assign Ycmow6 = (Ipfow6 | Bb0iu6);
assign Rcmow6 = (Rqfow6 | Ib0iu6);
assign Bbmow6 = (~(HRDATA[10] & Q2eow6));
assign Z2mow6 = (Fdmow6 & Dldow6);
assign Dldow6 = (~(H5how6 & Mdmow6));
assign Mdmow6 = (~(Tdmow6 & C6how6));
assign C6how6 = (~(Aemow6 & V3xhu6));
assign Aemow6 = (Hemow6 & Ktcow6);
assign Tdmow6 = (~(Oemow6 & Vemow6));
assign Vemow6 = (Cfmow6 & Dahow6);
assign Cfmow6 = (Tzlow6 & K3how6);
assign Tzlow6 = (Ny3ju6 | Ktcow6);
assign Ny3ju6 = (Fg3ju6 | R3how6);
assign Fg3ju6 = (~(Jfmow6 & Ej3ju6));
assign Oemow6 = (Qfmow6 & O1low6);
assign Qfmow6 = (~(Xfmow6 & Ktcow6));
assign Xfmow6 = (Egmow6 & Lgmow6);
assign Lgmow6 = (~(Sgmow6 & C0ehu6));
assign Sgmow6 = (~(Mjfiu6 | Cyfpw6[0]));
assign Egmow6 = (Rn2ju6 | Tfjiu6);
assign H5how6 = (~(Zgmow6 & Ghmow6));
assign Ghmow6 = (Nhmow6 & Uhmow6);
assign Uhmow6 = (Bimow6 | Q88ow6);
assign Q88ow6 = (Iimow6 & Pimow6);
assign Pimow6 = (Iydow6 | Ggtiu6);
assign Ggtiu6 = (Wimow6 & Djmow6);
assign Djmow6 = (Kjmow6 & Rjmow6);
assign Rjmow6 = (Yjmow6 & Fkmow6);
assign Fkmow6 = (Mkmow6 & Tkmow6);
assign Tkmow6 = (~(E1fiu6 & R4gpw6[43]));
assign Mkmow6 = (~(Q0fiu6 & R4gpw6[51]));
assign Yjmow6 = (Almow6 & Hlmow6);
assign Hlmow6 = (~(Tzdiu6 & R4gpw6[3]));
assign Almow6 = (~(STCALIB[15] & H1eow6));
assign Kjmow6 = (Olmow6 & Vlmow6);
assign Vlmow6 = (Cmmow6 & Jmmow6);
assign Jmmow6 = (P6ciu6 | Qkgiu6);
assign P6ciu6 = (~(Ydeow6 & Qmmow6));
assign Qmmow6 = (~(Xmmow6 & J1fow6));
assign J1fow6 = (!Feeow6);
assign Feeow6 = (~(O8low6 & A8low6));
assign Xmmow6 = (Meeow6 ? H7fow6 : B4fow6);
assign Ydeow6 = (A0fow6 & V0fow6);
assign A0fow6 = (~(Righu6 | Ahghu6));
assign Cmmow6 = (~(I3fiu6 & R4gpw6[11]));
assign Olmow6 = (Enmow6 & Lnmow6);
assign Lnmow6 = (~(G2fiu6 & R4gpw6[27]));
assign Enmow6 = (~(U2fiu6 & R4gpw6[19]));
assign Wimow6 = (Snmow6 & Znmow6);
assign Znmow6 = (Gomow6 & Nomow6);
assign Nomow6 = (Uomow6 & Bpmow6);
assign Bpmow6 = (~(Odgpw6[15] & M0eow6));
assign Uomow6 = (~(Tzfpw6[15] & Yvgiu6));
assign Gomow6 = (Ipmow6 & Ppmow6);
assign Ppmow6 = (~(F0eow6 & Vbgpw6[15]));
assign Ipmow6 = (~(Bagpw6[15] & M6eiu6));
assign Snmow6 = (Wpmow6 & Dqmow6);
assign Dqmow6 = (Kqmow6 & Rqmow6);
assign Rqmow6 = (~(C0fiu6 & R4gpw6[59]));
assign Kqmow6 = (~(Zlghu6 & Xrgiu6));
assign Xrgiu6 = (Yqmow6 & Ynhiu6);
assign Yqmow6 = (K5eiu6 & Jfgpw6[4]);
assign Wpmow6 = (Qgeow6 & Frmow6);
assign Frmow6 = (~(S1fiu6 & R4gpw6[35]));
assign Iimow6 = (Mrmow6 & Trmow6);
assign Trmow6 = (We3ju6 | Hfeow6);
assign We3ju6 = (!Y83ju6);
assign Y83ju6 = (Hv3ju6 ? L44ju6 : Re4ju6);
assign L44ju6 = (~(Asmow6 & Hsmow6));
assign Hsmow6 = (Osmow6 & Vsmow6);
assign Vsmow6 = (Ipfow6 | J80iu6);
assign Osmow6 = (Rqfow6 | Q80iu6);
assign Asmow6 = (Ctmow6 & Jtmow6);
assign Jtmow6 = (Ppfow6 | L90iu6);
assign Ctmow6 = (Kqfow6 | X80iu6);
assign Re4ju6 = (~(Qtmow6 & Xtmow6));
assign Xtmow6 = (Eumow6 & Lumow6);
assign Lumow6 = (Ipfow6 | S90iu6);
assign Eumow6 = (Rqfow6 | Z90iu6);
assign Qtmow6 = (Sumow6 & Zumow6);
assign Zumow6 = (Ppfow6 | Na0iu6);
assign Sumow6 = (Kqfow6 | Ga0iu6);
assign Mrmow6 = (~(Q2eow6 & HRDATA[15]));
assign Bimow6 = (Gvmow6 & Nvmow6);
assign Nvmow6 = (~(S2ziu6 & Cyfpw6[3]));
assign S2ziu6 = (~(Tfjiu6 | Hs0iu6));
assign Gvmow6 = (~(Uvmow6 & Yahow6));
assign Nhmow6 = (Bwmow6 & Bz3ju6);
assign Bwmow6 = (~(Iwmow6 & X88ow6));
assign X88ow6 = (~(Pwmow6 & Wwmow6));
assign Wwmow6 = (Iydow6 | Pxriu6);
assign Pxriu6 = (Dxmow6 & Kxmow6);
assign Kxmow6 = (Rxmow6 & Yxmow6);
assign Yxmow6 = (Fymow6 & Mymow6);
assign Mymow6 = (Tymow6 & Azmow6);
assign Azmow6 = (~(Odgpw6[7] & M0eow6));
assign Tymow6 = (~(Q0fiu6 & R4gpw6[49]));
assign Fymow6 = (Hzmow6 & Ozmow6);
assign Ozmow6 = (~(Bagpw6[7] & M6eiu6));
assign Hzmow6 = (~(C0fiu6 & R4gpw6[57]));
assign Rxmow6 = (Vzmow6 & C0now6);
assign C0now6 = (~(E1fiu6 & R4gpw6[41]));
assign Vzmow6 = (J0now6 & Q0now6);
assign Q0now6 = (~(Tzfpw6[7] & Yvgiu6));
assign J0now6 = (~(STCALIB[7] & H1eow6));
assign Dxmow6 = (X0now6 & E1now6);
assign E1now6 = (L1now6 & S1now6);
assign S1now6 = (~(F0eow6 & Vbgpw6[7]));
assign L1now6 = (Z1now6 & G2now6);
assign G2now6 = (~(S1fiu6 & R4gpw6[33]));
assign Z1now6 = (~(G2fiu6 & R4gpw6[25]));
assign X0now6 = (N2now6 & U2now6);
assign U2now6 = (~(U2fiu6 & R4gpw6[17]));
assign N2now6 = (B3now6 & I3now6);
assign I3now6 = (~(I3fiu6 & R4gpw6[9]));
assign B3now6 = (~(Tzdiu6 & R4gpw6[1]));
assign Pwmow6 = (P3now6 & W3now6);
assign W3now6 = (~(C2eow6 & Jb3ju6));
assign Jb3ju6 = (Hv3ju6 ? Ag4ju6 : Jw3ju6);
assign Ag4ju6 = (~(D4now6 & K4now6));
assign K4now6 = (R4now6 & Y4now6);
assign Y4now6 = (Ppfow6 | Pb0iu6);
assign Pb0iu6 = (F5now6 & M5now6);
assign M5now6 = (T5now6 & A6now6);
assign A6now6 = (H6now6 & O6now6);
assign O6now6 = (~(V6now6 & vis_r2_o[11]));
assign H6now6 = (~(C7now6 & vis_r6_o[11]));
assign T5now6 = (J7now6 & Q7now6);
assign Q7now6 = (~(X7now6 & vis_r5_o[11]));
assign J7now6 = (~(E8now6 & vis_r4_o[11]));
assign F5now6 = (L8now6 & S8now6);
assign S8now6 = (Z8now6 & G9now6);
assign G9now6 = (~(N9now6 & vis_r1_o[11]));
assign Z8now6 = (~(U9now6 & vis_r0_o[11]));
assign L8now6 = (Banow6 & Ianow6);
assign Ianow6 = (~(Panow6 & vis_r3_o[11]));
assign Banow6 = (~(Wanow6 & vis_r7_o[11]));
assign R4now6 = (Ipfow6 | Ua0iu6);
assign D4now6 = (Dbnow6 & Kbnow6);
assign Kbnow6 = (Rqfow6 | Bb0iu6);
assign Dbnow6 = (Kqfow6 | Ib0iu6);
assign Jw3ju6 = (~(Rbnow6 & Ybnow6));
assign Ybnow6 = (Fcnow6 & Mcnow6);
assign Mcnow6 = (Ppfow6 | I40iu6);
assign Fcnow6 = (Kqfow6 | B40iu6);
assign Rbnow6 = (Tcnow6 & Adnow6);
assign Adnow6 = (Ipfow6 | Wb0iu6);
assign Wb0iu6 = (Hdnow6 & Odnow6);
assign Odnow6 = (Vdnow6 & Cenow6);
assign Cenow6 = (Jenow6 & Qenow6);
assign Qenow6 = (~(V6now6 & vis_r2_o[10]));
assign Jenow6 = (~(C7now6 & vis_r6_o[10]));
assign Vdnow6 = (Xenow6 & Efnow6);
assign Efnow6 = (~(X7now6 & vis_r5_o[10]));
assign Xenow6 = (~(E8now6 & vis_r4_o[10]));
assign Hdnow6 = (Lfnow6 & Sfnow6);
assign Sfnow6 = (Zfnow6 & Ggnow6);
assign Ggnow6 = (~(N9now6 & vis_r1_o[10]));
assign Zfnow6 = (~(U9now6 & vis_r0_o[10]));
assign Lfnow6 = (Ngnow6 & Ugnow6);
assign Ugnow6 = (~(Panow6 & vis_r3_o[10]));
assign Ngnow6 = (~(Wanow6 & vis_r7_o[10]));
assign Tcnow6 = (Rqfow6 | U30iu6);
assign P3now6 = (~(HRDATA[7] & Q2eow6));
assign Iwmow6 = (~(Rn2ju6 & Bhnow6));
assign Bhnow6 = (~(Ihnow6 & Tfjiu6));
assign Ihnow6 = (~(Tr0iu6 & Phnow6));
assign Phnow6 = (Iwfpw6[0] | Iwfpw6[1]);
assign Rn2ju6 = (!A3aju6);
assign Zgmow6 = (Whnow6 & Dinow6);
assign Dinow6 = (~(Iwfpw6[1] & Kinow6));
assign Kinow6 = (~(Rinow6 & Yinow6));
assign Yinow6 = (~(Fjnow6 & Qyniu6));
assign Fjnow6 = (~(H78ow6 | Iwfpw6[0]));
assign H78ow6 = (Mjnow6 & Tjnow6);
assign Tjnow6 = (Iydow6 | N0viu6);
assign N0viu6 = (Aknow6 & Hknow6);
assign Hknow6 = (Oknow6 & Vknow6);
assign Vknow6 = (Clnow6 & Jlnow6);
assign Jlnow6 = (Qlnow6 & Xlnow6);
assign Xlnow6 = (~(Odgpw6[23] & M0eow6));
assign Qlnow6 = (~(Q0fiu6 & R4gpw6[53]));
assign Clnow6 = (Emnow6 & Lmnow6);
assign Lmnow6 = (~(Tzdiu6 & R4gpw6[5]));
assign Emnow6 = (~(I3fiu6 & R4gpw6[13]));
assign Oknow6 = (Smnow6 & Zmnow6);
assign Zmnow6 = (Gnnow6 & Nnnow6);
assign Nnnow6 = (~(Hqgiu6 & L1gpw6[1]));
assign Gnnow6 = (~(STCALIB[23] & H1eow6));
assign Smnow6 = (Unnow6 & Bonow6);
assign Bonow6 = (~(G2fiu6 & R4gpw6[29]));
assign Unnow6 = (~(U2fiu6 & R4gpw6[21]));
assign Aknow6 = (Ionow6 & Ponow6);
assign Ponow6 = (Wonow6 & Dpnow6);
assign Dpnow6 = (Kpnow6 & Rpnow6);
assign Rpnow6 = (~(Tzfpw6[23] & Yvgiu6));
assign Kpnow6 = (Qkgiu6 | U6piu6);
assign Wonow6 = (Ypnow6 & Fqnow6);
assign Fqnow6 = (~(Bagpw6[23] & M6eiu6));
assign Ypnow6 = (~(E1fiu6 & R4gpw6[45]));
assign Ionow6 = (Mqnow6 & Tqnow6);
assign Tqnow6 = (~(S1fiu6 & R4gpw6[37]));
assign Mqnow6 = (Arnow6 & Hrnow6);
assign Hrnow6 = (~(C0fiu6 & R4gpw6[61]));
assign Arnow6 = (~(F0eow6 & Vbgpw6[23]));
assign Mjnow6 = (Ornow6 & Vrnow6);
assign Vrnow6 = (Hfeow6 | Ha3ju6);
assign Ha3ju6 = (Hv3ju6 ? Csnow6 : C34ju6);
assign Csnow6 = (Ecjow6 & Lcjow6);
assign Lcjow6 = (Jsnow6 & Qsnow6);
assign Qsnow6 = (Ipfow6 | Y50iu6);
assign Jsnow6 = (Rqfow6 | M60iu6);
assign Ecjow6 = (Xsnow6 & Etnow6);
assign Etnow6 = (Ppfow6 | A70iu6);
assign Xsnow6 = (~(C3kow6 & Ltnow6));
assign C34ju6 = (Stnow6 & Ztnow6);
assign Ztnow6 = (Gunow6 & Nunow6);
assign Nunow6 = (Ipfow6 | H70iu6);
assign Gunow6 = (Rqfow6 | O70iu6);
assign Stnow6 = (Uunow6 & Bvnow6);
assign Bvnow6 = (Ppfow6 | C80iu6);
assign Uunow6 = (Kqfow6 | V70iu6);
assign Ornow6 = (~(HRDATA[23] & Q2eow6));
assign Rinow6 = (~(Uvmow6 & V78ow6));
assign V78ow6 = (~(Ivnow6 & Pvnow6));
assign Pvnow6 = (Iydow6 | Rw1iu6);
assign Rw1iu6 = (Wvnow6 & Dwnow6);
assign Dwnow6 = (Kwnow6 & Rwnow6);
assign Rwnow6 = (Ywnow6 & Fxnow6);
assign Fxnow6 = (Mxnow6 & Txnow6);
assign Txnow6 = (Te6iu6 | Qkgiu6);
assign Mxnow6 = (~(Hqgiu6 & H8gpw6[1]));
assign Hqgiu6 = (Aynow6 & Ynhiu6);
assign Aynow6 = (K5eiu6 & U89iu6);
assign Ywnow6 = (Hynow6 & Oynow6);
assign Oynow6 = (~(STCALIB[25] & H1eow6));
assign Hynow6 = (~(C0fiu6 & R4gpw6[63]));
assign C0fiu6 = (Vynow6 & Cznow6);
assign Kwnow6 = (Jznow6 & Qznow6);
assign Qznow6 = (~(S1fiu6 & R4gpw6[39]));
assign S1fiu6 = (Xznow6 & Vynow6);
assign Jznow6 = (E0oow6 & L0oow6);
assign L0oow6 = (~(Tzdiu6 & R4gpw6[7]));
assign Tzdiu6 = (Xznow6 & Pjyiu6);
assign E0oow6 = (~(Q0fiu6 & R4gpw6[55]));
assign Q0fiu6 = (S0oow6 & Vynow6);
assign Wvnow6 = (Z0oow6 & G1oow6);
assign G1oow6 = (N1oow6 & U1oow6);
assign U1oow6 = (B2oow6 & I2oow6);
assign I2oow6 = (~(Pceow6 & P2oow6));
assign P2oow6 = (Nzhiu6 | Vbgpw6[31]);
assign B2oow6 = (~(G2fiu6 & R4gpw6[31]));
assign G2fiu6 = (Pjyiu6 & Cznow6);
assign N1oow6 = (W2oow6 & D3oow6);
assign D3oow6 = (~(U2fiu6 & R4gpw6[23]));
assign U2fiu6 = (S0oow6 & Pjyiu6);
assign S0oow6 = (K3oow6 & Jfgpw6[3]);
assign K3oow6 = (~(Jfgpw6[2] | Jfgpw6[4]));
assign W2oow6 = (~(E1fiu6 & R4gpw6[47]));
assign E1fiu6 = (Vynow6 & Dtjow6);
assign Z0oow6 = (R3oow6 & Y3oow6);
assign Y3oow6 = (Tpgiu6 | F4oow6);
assign Tpgiu6 = (~(Rzciu6 & Cznow6));
assign R3oow6 = (M4oow6 & T4oow6);
assign T4oow6 = (~(I3fiu6 & R4gpw6[15]));
assign I3fiu6 = (Pjyiu6 & Dtjow6);
assign M4oow6 = (~(Odgpw6[31] & M0eow6));
assign Ivnow6 = (A5oow6 & H5oow6);
assign H5oow6 = (Hfeow6 | Mg3ju6);
assign Mg3ju6 = (!O5oow6);
assign O5oow6 = (V5oow6 ? Vh3ju6 : Qb3ju6);
assign V5oow6 = (Queow6 & Solow6);
assign Solow6 = (~(V2kow6 & Ppfow6));
assign Queow6 = (C6oow6 & Cyfpw6[3]);
assign C6oow6 = (J6oow6 & Hzfow6);
assign J6oow6 = (Azfow6 | Ppfow6);
assign Vh3ju6 = (!Bz3ju6);
assign Qb3ju6 = (Hv3ju6 ? Lx3ju6 : Vajow6);
assign Lx3ju6 = (~(Q6oow6 & X6oow6));
assign X6oow6 = (E7oow6 & L7oow6);
assign L7oow6 = (Rqfow6 | W40iu6);
assign E7oow6 = (Kqfow6 | D50iu6);
assign Q6oow6 = (S7oow6 & Z7oow6);
assign Z7oow6 = (Ppfow6 | K50iu6);
assign S7oow6 = (Ipfow6 | P40iu6);
assign Vajow6 = (~(G8oow6 & N8oow6));
assign N8oow6 = (U8oow6 & B9oow6);
assign B9oow6 = (Ipfow6 | F60iu6);
assign U8oow6 = (Rqfow6 | E90iu6);
assign G8oow6 = (I9oow6 & P9oow6);
assign P9oow6 = (Ppfow6 | R50iu6);
assign I9oow6 = (Kqfow6 | Dc0iu6);
assign A5oow6 = (~(Q2eow6 & HRDATA[31]));
assign Uvmow6 = (~(W9oow6 & Daoow6));
assign Daoow6 = (X5oiu6 | Cyfpw6[0]);
assign W9oow6 = (~(Iwfpw6[0] & Qyniu6));
assign Whnow6 = (~(V3xhu6 & Hemow6));
assign Fdmow6 = (Gkcow6 | Uqdow6);
assign Uqdow6 = (!Mmdow6);
assign Mmdow6 = (~(Hlziu6 & Rahow6));
assign Rahow6 = (~(Kaoow6 & Ktcow6));
assign Kaoow6 = (Fd0iu6 & Pthiu6);
assign Hlziu6 = (O1low6 & W9how6);
assign W9how6 = (~(Ktcow6 & Vxniu6));
assign O1low6 = (Kf3ju6 | Ktcow6);
assign Kf3ju6 = (X6how6 | Df3ju6);
assign X6how6 = (~(Raoow6 & Oa3ju6));
assign Raoow6 = (F93ju6 & U54ju6);
assign Gkcow6 = (Yaoow6 & Fboow6);
assign Fboow6 = (Mboow6 & Tboow6);
assign Tboow6 = (Rcfow6 | Yt3ju6);
assign Yt3ju6 = (Acoow6 & Hcoow6);
assign Hcoow6 = (Ocoow6 & Vcoow6);
assign Vcoow6 = (Kqfow6 | I40iu6);
assign I40iu6 = (Cdoow6 & Jdoow6);
assign Jdoow6 = (Qdoow6 & Xdoow6);
assign Xdoow6 = (Eeoow6 & Leoow6);
assign Leoow6 = (~(V6now6 & vis_r2_o[7]));
assign Eeoow6 = (~(C7now6 & vis_r6_o[7]));
assign Qdoow6 = (Seoow6 & Zeoow6);
assign Zeoow6 = (~(X7now6 & vis_r5_o[7]));
assign Seoow6 = (~(E8now6 & vis_r4_o[7]));
assign Cdoow6 = (Gfoow6 & Nfoow6);
assign Nfoow6 = (Ufoow6 & Bgoow6);
assign Bgoow6 = (~(N9now6 & vis_r1_o[7]));
assign Ufoow6 = (~(U9now6 & vis_r0_o[7]));
assign Gfoow6 = (Igoow6 & Pgoow6);
assign Pgoow6 = (~(Panow6 & vis_r3_o[7]));
assign Igoow6 = (~(Wanow6 & vis_r7_o[7]));
assign Ocoow6 = (Rqfow6 | B40iu6);
assign B40iu6 = (Wgoow6 & Dhoow6);
assign Dhoow6 = (Khoow6 & Rhoow6);
assign Rhoow6 = (Yhoow6 & Fioow6);
assign Fioow6 = (~(V6now6 & vis_r2_o[8]));
assign Yhoow6 = (~(C7now6 & vis_r6_o[8]));
assign Khoow6 = (Mioow6 & Tioow6);
assign Tioow6 = (~(X7now6 & vis_r5_o[8]));
assign Mioow6 = (~(E8now6 & vis_r4_o[8]));
assign Wgoow6 = (Ajoow6 & Hjoow6);
assign Hjoow6 = (Ojoow6 & Vjoow6);
assign Vjoow6 = (~(N9now6 & vis_r1_o[8]));
assign Ojoow6 = (~(U9now6 & vis_r0_o[8]));
assign Ajoow6 = (Ckoow6 & Jkoow6);
assign Jkoow6 = (~(Panow6 & vis_r3_o[8]));
assign Ckoow6 = (~(Wanow6 & vis_r7_o[8]));
assign Acoow6 = (Qkoow6 & Xkoow6);
assign Xkoow6 = (Ipfow6 | U30iu6);
assign Qkoow6 = (Ppfow6 | P40iu6);
assign Mboow6 = (Iydow6 | Jaqiu6);
assign Jaqiu6 = (Eloow6 & Lloow6);
assign Lloow6 = (Sloow6 & Zloow6);
assign Zloow6 = (Gmoow6 & Nmoow6);
assign Nmoow6 = (~(Odgpw6[2] & M0eow6));
assign Gmoow6 = (Umoow6 & Bnoow6);
assign Bnoow6 = (~(Ndghu6 & Fpgiu6));
assign Fpgiu6 = (Rzciu6 & Xznow6);
assign Umoow6 = (~(STCALIB[2] & H1eow6));
assign Sloow6 = (Inoow6 & Pnoow6);
assign Pnoow6 = (~(ECOREVNUM[2] & I5eow6));
assign Inoow6 = (~(Y5eiu6 & Wnoow6));
assign Wnoow6 = (STCALIB[25] | Ftghu6);
assign Y5eiu6 = (Vynow6 & Wjyiu6);
assign Eloow6 = (Dooow6 & Kooow6);
assign Kooow6 = (Rooow6 & Yooow6);
assign Yooow6 = (~(F0eow6 & Vbgpw6[2]));
assign Rooow6 = (~(Bagpw6[2] & M6eiu6));
assign Dooow6 = (Fpoow6 & Mpoow6);
assign Mpoow6 = (~(Tzfpw6[2] & Yvgiu6));
assign Fpoow6 = (Qkgiu6 | Tfciu6);
assign Yaoow6 = (Tpoow6 & Aqoow6);
assign Aqoow6 = (~(Qtfow6 & Zx3ju6));
assign Zx3ju6 = (~(Hqoow6 & Oqoow6));
assign Oqoow6 = (Vqoow6 & Croow6);
assign Croow6 = (Ipfow6 | W40iu6);
assign W40iu6 = (Jroow6 & Qroow6);
assign Qroow6 = (Xroow6 & Esoow6);
assign Esoow6 = (Lsoow6 & Ssoow6);
assign Ssoow6 = (~(V6now6 & vis_r2_o[5]));
assign Lsoow6 = (~(C7now6 & vis_r6_o[5]));
assign Xroow6 = (Zsoow6 & Gtoow6);
assign Gtoow6 = (~(X7now6 & vis_r5_o[5]));
assign Zsoow6 = (~(E8now6 & vis_r4_o[5]));
assign Jroow6 = (Ntoow6 & Utoow6);
assign Utoow6 = (Buoow6 & Iuoow6);
assign Iuoow6 = (~(N9now6 & vis_r1_o[5]));
assign Buoow6 = (~(U9now6 & vis_r0_o[5]));
assign Ntoow6 = (Puoow6 & Wuoow6);
assign Wuoow6 = (~(Panow6 & vis_r3_o[5]));
assign Puoow6 = (~(Wanow6 & vis_r7_o[5]));
assign Vqoow6 = (Kqfow6 | K50iu6);
assign K50iu6 = (Dvoow6 & Kvoow6);
assign Kvoow6 = (Rvoow6 & Yvoow6);
assign Yvoow6 = (Fwoow6 & Mwoow6);
assign Mwoow6 = (~(V6now6 & vis_r2_o[3]));
assign Fwoow6 = (~(C7now6 & vis_r6_o[3]));
assign Rvoow6 = (Twoow6 & Axoow6);
assign Axoow6 = (~(X7now6 & vis_r5_o[3]));
assign Twoow6 = (~(E8now6 & vis_r4_o[3]));
assign Dvoow6 = (Hxoow6 & Oxoow6);
assign Oxoow6 = (Vxoow6 & Cyoow6);
assign Cyoow6 = (~(N9now6 & vis_r1_o[3]));
assign Vxoow6 = (~(U9now6 & vis_r0_o[3]));
assign Hxoow6 = (Jyoow6 & Qyoow6);
assign Qyoow6 = (~(Panow6 & vis_r3_o[3]));
assign Jyoow6 = (~(Wanow6 & vis_r7_o[3]));
assign Hqoow6 = (Xyoow6 & Ezoow6);
assign Ezoow6 = (Ppfow6 | F60iu6);
assign F60iu6 = (Lzoow6 & Szoow6);
assign Szoow6 = (Zzoow6 & G0pow6);
assign G0pow6 = (N0pow6 & U0pow6);
assign U0pow6 = (~(V6now6 & vis_r2_o[2]));
assign N0pow6 = (~(C7now6 & vis_r6_o[2]));
assign Zzoow6 = (B1pow6 & I1pow6);
assign I1pow6 = (~(X7now6 & vis_r5_o[2]));
assign B1pow6 = (~(E8now6 & vis_r4_o[2]));
assign Lzoow6 = (P1pow6 & W1pow6);
assign W1pow6 = (D2pow6 & K2pow6);
assign K2pow6 = (~(N9now6 & vis_r1_o[2]));
assign D2pow6 = (~(U9now6 & vis_r0_o[2]));
assign P1pow6 = (R2pow6 & Y2pow6);
assign Y2pow6 = (~(Panow6 & vis_r3_o[2]));
assign R2pow6 = (~(Wanow6 & vis_r7_o[2]));
assign Xyoow6 = (Rqfow6 | D50iu6);
assign D50iu6 = (F3pow6 & M3pow6);
assign M3pow6 = (T3pow6 & A4pow6);
assign A4pow6 = (H4pow6 & O4pow6);
assign O4pow6 = (~(V6now6 & vis_r2_o[4]));
assign H4pow6 = (~(C7now6 & vis_r6_o[4]));
assign T3pow6 = (V4pow6 & C5pow6);
assign C5pow6 = (~(X7now6 & vis_r5_o[4]));
assign V4pow6 = (~(E8now6 & vis_r4_o[4]));
assign F3pow6 = (J5pow6 & Q5pow6);
assign Q5pow6 = (X5pow6 & E6pow6);
assign E6pow6 = (~(N9now6 & vis_r1_o[4]));
assign X5pow6 = (~(U9now6 & vis_r0_o[4]));
assign J5pow6 = (L6pow6 & S6pow6);
assign S6pow6 = (~(Panow6 & vis_r3_o[4]));
assign L6pow6 = (~(Wanow6 & vis_r7_o[4]));
assign Tpoow6 = (~(HRDATA[2] & Q2eow6));
assign L2mow6 = (Z6pow6 & G7pow6);
assign G7pow6 = (Wlcow6 | Kldow6);
assign Kldow6 = (Dtcow6 & Dahow6);
assign Dahow6 = (Ch4ju6 | Ktcow6);
assign Ch4ju6 = (Avcow6 | R3how6);
assign R3how6 = (~(Mr0iu6 | N7pow6));
assign Avcow6 = (~(Jfmow6 & F93ju6));
assign Jfmow6 = (M93ju6 & U54ju6);
assign M93ju6 = (!Oa3ju6);
assign Dtcow6 = (Tucow6 | Qxaiu6);
assign Wlcow6 = (U7pow6 & B8pow6);
assign B8pow6 = (I8pow6 & P8pow6);
assign P8pow6 = (Rcfow6 | R04ju6);
assign R04ju6 = (W8pow6 & D9pow6);
assign D9pow6 = (K9pow6 & R9pow6);
assign R9pow6 = (Ipfow6 | O70iu6);
assign K9pow6 = (Rqfow6 | V70iu6);
assign W8pow6 = (Y9pow6 & Fapow6);
assign Fapow6 = (Ppfow6 | J80iu6);
assign Y9pow6 = (Kqfow6 | C80iu6);
assign Rcfow6 = (!Dyeow6);
assign Dyeow6 = (~(Hfeow6 | J2eow6));
assign I8pow6 = (Iydow6 | U1uiu6);
assign U1uiu6 = (Mapow6 & Tapow6);
assign Tapow6 = (Abpow6 & Hbpow6);
assign Hbpow6 = (~(Pceow6 & Obpow6));
assign Obpow6 = (Nzhiu6 | Vbgpw6[18]);
assign Pceow6 = (Nzhiu6 | F0eow6);
assign Abpow6 = (Vbpow6 & Ccpow6);
assign Ccpow6 = (~(Tzfpw6[18] & Yvgiu6));
assign Yvgiu6 = (Jcpow6 & Vynow6);
assign Jcpow6 = (Ynhiu6 & U89iu6);
assign Vbpow6 = (~(Odgpw6[18] & M0eow6));
assign Mapow6 = (Qcpow6 & Qgeow6);
assign Qgeow6 = (!I5eow6);
assign I5eow6 = (~(Xcpow6 & Edpow6));
assign Edpow6 = (~(Ldpow6 & Cpwiu6));
assign Cpwiu6 = (Sdpow6 & X8hpw6[5]);
assign Sdpow6 = (~(X8hpw6[0] | X8hpw6[6]));
assign Ldpow6 = (Ilwiu6 & Q4wiu6);
assign Q4wiu6 = (~(X8hpw6[1] | X8hpw6[4]));
assign Ilwiu6 = (X8hpw6[2] & Vm6iu6);
assign Vm6iu6 = (!X8hpw6[3]);
assign Xcpow6 = (~(Xznow6 & K5eiu6));
assign Xznow6 = (Zdpow6 & Jfgpw6[2]);
assign Qcpow6 = (Gepow6 & Nepow6);
assign Nepow6 = (~(Bagpw6[18] & M6eiu6));
assign M6eiu6 = (Vynow6 & D5eiu6);
assign Gepow6 = (~(STCALIB[18] & H1eow6));
assign H1eow6 = (Uepow6 & Vynow6);
assign Vynow6 = (~(Uh7iu6 | Jfgpw6[1]));
assign Uepow6 = (Ynhiu6 & Jfgpw6[4]);
assign Ynhiu6 = (Jfgpw6[3] & Jfgpw6[2]);
assign U7pow6 = (Bfpow6 & Ifpow6);
assign Ifpow6 = (~(Qtfow6 & Ye4ju6));
assign Ye4ju6 = (~(Pfpow6 & Wfpow6));
assign Wfpow6 = (Dgpow6 & Kgpow6);
assign Kgpow6 = (Ipfow6 | Q80iu6);
assign Dgpow6 = (Ppfow6 | S90iu6);
assign Pfpow6 = (Rgpow6 & Ygpow6);
assign Ygpow6 = (Kqfow6 | L90iu6);
assign Rgpow6 = (Rqfow6 | X80iu6);
assign Qtfow6 = (~(Hfeow6 | Hv3ju6));
assign Hfeow6 = (!C2eow6);
assign Bfpow6 = (~(HRDATA[18] & Q2eow6));
assign Z6pow6 = (Ukcow6 | Spdow6);
assign Spdow6 = (!Fmdow6);
assign Fmdow6 = (~(Fhpow6 & Mhpow6));
assign Mhpow6 = (~(T4how6 & Cyfpw6[3]));
assign T4how6 = (Thpow6 & Iwfpw6[1]);
assign Thpow6 = (~(Tucow6 | Cyfpw6[1]));
assign Fhpow6 = (F4how6 & K3how6);
assign K3how6 = (L7how6 | Ktcow6);
assign Ktcow6 = (!Tucow6);
assign L7how6 = (!Pe3ju6);
assign Pe3ju6 = (Aipow6 & Oa3ju6);
assign Aipow6 = (Ej3ju6 & U54ju6);
assign U54ju6 = (Ii0iu6 | Z53ju6);
assign Z53ju6 = (!Q43ju6);
assign Q43ju6 = (~(Hipow6 & Oipow6));
assign Oipow6 = (~(Vipow6 & Cjpow6));
assign Cjpow6 = (Jjpow6 & Qjpow6);
assign Qjpow6 = (~(S8fpw6[4] | H4ghu6));
assign Jjpow6 = (~(S8fpw6[2] | S8fpw6[3]));
assign Vipow6 = (Xjpow6 & Pugiu6);
assign Xjpow6 = (~(S8fpw6[0] | S8fpw6[1]));
assign Hipow6 = (Ekpow6 & Zc3ju6);
assign Zc3ju6 = (~(Pfoiu6 & Lkpow6));
assign Lkpow6 = (~(Zvzhu6 & Svzhu6));
assign Ekpow6 = (Yn2ju6 | Gwzhu6);
assign F4how6 = (~(Skpow6 & Zkpow6));
assign Zkpow6 = (~(Wmaiu6 | Tr0iu6));
assign Wmaiu6 = (!Glpow6);
assign Skpow6 = (~(Yahow6 | Tucow6));
assign Tucow6 = (~(Qcoiu6 & Nlpow6));
assign Nlpow6 = (~(Ulpow6 & Xkaow6));
assign Ulpow6 = (~(Imaiu6 | Y7ghu6));
assign Qcoiu6 = (!Bmpow6);
assign Yahow6 = (!Iwfpw6[1]);
assign Ukcow6 = (Impow6 & Pmpow6);
assign Pmpow6 = (Iydow6 | Wmviu6);
assign Wmviu6 = (Wmpow6 & Dnpow6);
assign Dnpow6 = (~(Odgpw6[26] & M0eow6));
assign M0eow6 = (Pjyiu6 & Knpow6);
assign Pjyiu6 = (Jfgpw6[0] & Jfgpw6[1]);
assign Wmpow6 = (Rnpow6 & Ynpow6);
assign Ynpow6 = (~(F0eow6 & Vbgpw6[26]));
assign F0eow6 = (K5eiu6 & Knpow6);
assign Knpow6 = (Wjyiu6 | D5eiu6);
assign D5eiu6 = (Fopow6 & Jfgpw6[4]);
assign Fopow6 = (~(Jfgpw6[2] | Jfgpw6[3]));
assign Rnpow6 = (~(Yyghu6 & T7eow6));
assign T7eow6 = (!Qkgiu6);
assign Qkgiu6 = (~(K5eiu6 & Dtjow6));
assign Dtjow6 = (Mopow6 & Jfgpw6[4]);
assign Mopow6 = (~(Ka9iu6 | Jfgpw6[3]));
assign Iydow6 = (~(Hemow6 & Topow6));
assign Topow6 = (~(Rzciu6 & Wjyiu6));
assign Impow6 = (Appow6 & Hppow6);
assign Hppow6 = (~(C2eow6 & Oppow6));
assign Oppow6 = (~(Vppow6 & Cqpow6));
assign Cqpow6 = (Jqpow6 | Bz3ju6);
assign Bz3ju6 = (~(Qqpow6 & E5ehu6));
assign Qqpow6 = (~(Xqpow6 | R50iu6));
assign Xqpow6 = (~(F3aiu6 | Pt2ju6));
assign Vppow6 = (~(F84ju6 & Erpow6));
assign Erpow6 = (O24ju6 | Hv3ju6);
assign O24ju6 = (~(Lrpow6 & Srpow6));
assign Srpow6 = (Zrpow6 & Gspow6);
assign Gspow6 = (Ipfow6 | M60iu6);
assign Zrpow6 = (Ppfow6 | H70iu6);
assign Lrpow6 = (Nspow6 & Uspow6);
assign Uspow6 = (Kqfow6 | A70iu6);
assign Nspow6 = (Rqfow6 | T60iu6);
assign F84ju6 = (Btpow6 & Jqpow6);
assign Jqpow6 = (~(Itpow6 & Jbjow6));
assign Jbjow6 = (Ptpow6 & Cyfpw6[3]);
assign Ptpow6 = (Wtpow6 & Azfow6);
assign Azfow6 = (!Lveow6);
assign Lveow6 = (J2eow6 & Uieow6);
assign Uieow6 = (!V2kow6);
assign Wtpow6 = (Ppfow6 | V2kow6);
assign Itpow6 = (Kqfow6 ? Qbjow6 : V2kow6);
assign Qbjow6 = (Hzfow6 | Dupow6);
assign Hzfow6 = (~(V2kow6 & Hv3ju6));
assign V2kow6 = (~(N7pow6 | Df3ju6));
assign Df3ju6 = (Vwaiu6 & Mr0iu6);
assign N7pow6 = (Kupow6 & Rupow6);
assign Rupow6 = (~(F93ju6 | Oa3ju6));
assign Oa3ju6 = (H4ghu6 ? Yupow6 : X43ju6);
assign Yupow6 = (~(G63ju6 ^ Sc3ju6));
assign Sc3ju6 = (!X43ju6);
assign X43ju6 = (~(Fvpow6 & Mvpow6));
assign Mvpow6 = (Yn2ju6 | Nwzhu6);
assign Fvpow6 = (A4oiu6 | Qjoiu6);
assign F93ju6 = (!Ej3ju6);
assign Ej3ju6 = (H4ghu6 ? Awpow6 : Tvpow6);
assign Awpow6 = (~(Hwpow6 & G63ju6));
assign G63ju6 = (Owpow6 | Vwpow6);
assign Hwpow6 = (~(Vwpow6 & Owpow6));
assign Tvpow6 = (!Owpow6);
assign Owpow6 = (~(Cxpow6 & Jxpow6));
assign Jxpow6 = (Yn2ju6 | Uwzhu6);
assign Cxpow6 = (Cajiu6 | A4oiu6);
assign Cajiu6 = (!S8fpw6[3]);
assign Kupow6 = (~(Hv3ju6 | Ppfow6));
assign Hv3ju6 = (!J2eow6);
assign Btpow6 = (Eolow6 | J2eow6);
assign J2eow6 = (H4ghu6 ? Xxpow6 : Qxpow6);
assign Xxpow6 = (~(Eypow6 & Vwpow6));
assign Vwpow6 = (Lypow6 | Sypow6);
assign Eypow6 = (~(Sypow6 & Lypow6));
assign Lypow6 = (!Qxpow6);
assign Qxpow6 = (Zypow6 & Gzpow6);
assign Gzpow6 = (Yn2ju6 | Pxzhu6);
assign Zypow6 = (B5kiu6 | A4oiu6);
assign Eolow6 = (~(Nzpow6 & Uzpow6));
assign Uzpow6 = (B0qow6 & I0qow6);
assign I0qow6 = (Ipfow6 | E90iu6);
assign Ipfow6 = (P0qow6 | W0qow6);
assign B0qow6 = (Rqfow6 | Dc0iu6);
assign Rqfow6 = (!Gweow6);
assign Gweow6 = (~(D1qow6 | P0qow6));
assign Nzpow6 = (K1qow6 & R1qow6);
assign R1qow6 = (Ppfow6 | Y50iu6);
assign Ppfow6 = (!Dupow6);
assign Dupow6 = (P0qow6 & W0qow6);
assign K1qow6 = (Kqfow6 | R50iu6);
assign Kqfow6 = (!C3kow6);
assign C3kow6 = (P0qow6 & D1qow6);
assign P0qow6 = (H4ghu6 ? F2qow6 : Y1qow6);
assign F2qow6 = (~(M2qow6 & Sypow6));
assign Sypow6 = (~(Y1qow6 & W0qow6));
assign M2qow6 = (W0qow6 | Y1qow6);
assign W0qow6 = (!D1qow6);
assign D1qow6 = (~(T2qow6 & A3qow6));
assign A3qow6 = (Yn2ju6 | N30iu6);
assign T2qow6 = (Je8iu6 | A4oiu6);
assign Je8iu6 = (!S8fpw6[0]);
assign Y1qow6 = (H3qow6 & O3qow6);
assign O3qow6 = (Yn2ju6 | O00iu6);
assign H3qow6 = (Y8biu6 | A4oiu6);
assign Y8biu6 = (!S8fpw6[1]);
assign C2eow6 = (E5ehu6 & V3qow6);
assign V3qow6 = (~(C4qow6 & J4qow6));
assign J4qow6 = (Tr0iu6 | Gwyiu6);
assign C4qow6 = (~(Bmpow6 | A3aju6));
assign Bmpow6 = (Hs0iu6 & K9aiu6);
assign Appow6 = (~(HRDATA[26] & Q2eow6));
assign Q2eow6 = (Ytwiu6 & Hemow6);
assign Hemow6 = (~(Nm1ju6 | Q4qow6));
assign Q4qow6 = (~(X4qow6 | E5qow6));
assign E5qow6 = (Cyfpw6[1] ? Glpow6 : L5qow6);
assign Glpow6 = (Gwyiu6 & Nlaiu6);
assign L5qow6 = (~(S5qow6 | Hs0iu6));
assign X4qow6 = (~(Z5qow6 & K9aiu6));
assign Z5qow6 = (Xkaow6 | C0ehu6);
assign Nm1ju6 = (!E5ehu6);
assign Ytwiu6 = (Rzciu6 & Wjyiu6);
assign Wjyiu6 = (Zdpow6 & Ka9iu6);
assign Ka9iu6 = (!Jfgpw6[2]);
assign Zdpow6 = (~(Jfgpw6[3] | Jfgpw6[4]));
assign Rzciu6 = (~(Jfgpw6[0] | Jfgpw6[1]));
assign Zgziu6 = (~(Jmziu6 | Gu8iu6));
assign A0mow6 = (G6qow6 & N6qow6);
assign N6qow6 = (~(Zsfpw6[9] & Cmziu6));
assign Cmziu6 = (~(Hr8iu6 | Jmziu6));
assign Hr8iu6 = (Et8iu6 | U6qow6);
assign G6qow6 = (~(vis_pc_o[9] & Jmziu6));
assign Jmziu6 = (~(HREADY & B7qow6));
assign Acohu6 = (~(I7qow6 & P7qow6));
assign P7qow6 = (~(Umhow6 & HRDATA[19]));
assign I7qow6 = (~(Hrfpw6[3] & Qqhiu6));
assign Tbohu6 = (~(W7qow6 & D8qow6));
assign D8qow6 = (~(Umhow6 & HRDATA[18]));
assign W7qow6 = (~(Hrfpw6[2] & Qqhiu6));
assign Mbohu6 = (~(K8qow6 & R8qow6));
assign R8qow6 = (~(Umhow6 & HRDATA[17]));
assign Umhow6 = (~(Wz4iu6 | Qqhiu6));
assign Wz4iu6 = (!Glhiu6);
assign Glhiu6 = (Vobiu6 & Hs7iu6);
assign K8qow6 = (~(Hrfpw6[1] & Qqhiu6));
assign Fbohu6 = (Qqhiu6 ? Hrfpw6[14] : Rw8iu6);
assign Qqhiu6 = (~(Dxfhu6 & HREADY));
assign Rw8iu6 = (~(Hs7iu6 & Y8qow6));
assign Y8qow6 = (~(HRDATA[30] & Vobiu6));
assign Vobiu6 = (~(F9qow6 | N19iu6));
assign N19iu6 = (!vis_tbit_o);
assign F9qow6 = (V3xhu6 | Yyfhu6);
assign V3xhu6 = (HRESP & Qaxiu6);
assign Hs7iu6 = (!Aghhu6);
assign Yaohu6 = (~(Kaohu6 & M9qow6));
assign M9qow6 = (~(T9qow6 & G3eiu6));
assign G3eiu6 = (Npdhu6 & HWDATA[2]);
assign T9qow6 = (Uzhiu6 & Nzhiu6);
assign Nzhiu6 = (!Yreow6);
assign Yreow6 = (~(Cznow6 & K5eiu6));
assign K5eiu6 = (Jfgpw6[1] & Uh7iu6);
assign Uh7iu6 = (!Jfgpw6[0]);
assign Cznow6 = (Aaqow6 & Jfgpw6[3]);
assign Aaqow6 = (~(U89iu6 | Jfgpw6[2]));
assign U89iu6 = (!Jfgpw6[4]);
assign Uzhiu6 = (Haqow6 & Oaqow6);
assign Oaqow6 = (Vaqow6 & Cbqow6);
assign Cbqow6 = (Jbqow6 & Qbqow6);
assign Qbqow6 = (~(HWDATA[29] | HWDATA[16]));
assign HWDATA[16] = (~(Xbqow6 & Ecqow6));
assign Ecqow6 = (~(Lcqow6 & L35ju6));
assign Xbqow6 = (Scqow6 & Zcqow6);
assign Zcqow6 = (~(Gdqow6 & Xc9ju6));
assign Xc9ju6 = (~(Ndqow6 & Udqow6));
assign Udqow6 = (Beqow6 & Ieqow6);
assign Ieqow6 = (Peqow6 & Weqow6);
assign Weqow6 = (~(Fkfpw6[16] & Dfqow6));
assign Peqow6 = (Kfqow6 & Rfqow6);
assign Rfqow6 = (~(vis_psp_o[14] & Yfqow6));
assign Kfqow6 = (~(vis_msp_o[14] & Fgqow6));
assign Beqow6 = (Mgqow6 & Tgqow6);
assign Tgqow6 = (~(vis_r14_o[16] & Ahqow6));
assign Mgqow6 = (~(vis_r12_o[16] & Hhqow6));
assign Ndqow6 = (Ohqow6 & Vhqow6);
assign Vhqow6 = (Ciqow6 & Jiqow6);
assign Jiqow6 = (~(vis_r9_o[16] & Qiqow6));
assign Ciqow6 = (Xiqow6 & Ejqow6);
assign Ejqow6 = (~(vis_r11_o[16] & Ljqow6));
assign Xiqow6 = (~(vis_r10_o[16] & Sjqow6));
assign Ohqow6 = (Q10iu6 & Zjqow6);
assign Zjqow6 = (~(vis_r8_o[16] & Gkqow6));
assign Q10iu6 = (Nkqow6 & Ukqow6);
assign Ukqow6 = (Blqow6 & Ilqow6);
assign Ilqow6 = (Plqow6 & Wlqow6);
assign Wlqow6 = (~(vis_r2_o[16] & Dmqow6));
assign Plqow6 = (~(vis_r6_o[16] & Kmqow6));
assign Blqow6 = (Rmqow6 & Ymqow6);
assign Ymqow6 = (~(vis_r5_o[16] & Fnqow6));
assign Rmqow6 = (~(vis_r4_o[16] & Mnqow6));
assign Nkqow6 = (Tnqow6 & Aoqow6);
assign Aoqow6 = (Hoqow6 & Ooqow6);
assign Ooqow6 = (~(vis_r1_o[16] & Voqow6));
assign Hoqow6 = (~(vis_r0_o[16] & Cpqow6));
assign Tnqow6 = (Jpqow6 & Qpqow6);
assign Qpqow6 = (~(vis_r3_o[16] & Xpqow6));
assign Jpqow6 = (~(vis_r7_o[16] & Eqqow6));
assign Scqow6 = (~(Z54iu6 & R0nhu6));
assign Z54iu6 = (Shhpw6[16] & Iqzhu6);
assign HWDATA[29] = (~(Lqqow6 & Sqqow6));
assign Sqqow6 = (Zqqow6 & Grqow6);
assign Grqow6 = (~(Gdqow6 & Wh8iu6));
assign Wh8iu6 = (~(Nrqow6 & Urqow6));
assign Urqow6 = (Bsqow6 & Isqow6);
assign Isqow6 = (Psqow6 & Wsqow6);
assign Wsqow6 = (~(vis_r11_o[29] & Ljqow6));
assign Psqow6 = (Dtqow6 & Ktqow6);
assign Ktqow6 = (~(vis_r9_o[29] & Qiqow6));
assign Dtqow6 = (~(Fkfpw6[29] & Dfqow6));
assign Bsqow6 = (Rtqow6 & Ytqow6);
assign Ytqow6 = (~(vis_r10_o[29] & Sjqow6));
assign Rtqow6 = (~(vis_psp_o[27] & Yfqow6));
assign Nrqow6 = (Fuqow6 & Muqow6);
assign Muqow6 = (Tuqow6 & Avqow6);
assign Avqow6 = (~(vis_r12_o[29] & Hhqow6));
assign Tuqow6 = (Hvqow6 & Ovqow6);
assign Ovqow6 = (~(vis_msp_o[27] & Fgqow6));
assign Hvqow6 = (~(vis_r14_o[29] & Ahqow6));
assign Fuqow6 = (Wxzhu6 & Vvqow6);
assign Vvqow6 = (~(vis_r8_o[29] & Gkqow6));
assign Wxzhu6 = (Cwqow6 & Jwqow6);
assign Jwqow6 = (Qwqow6 & Xwqow6);
assign Xwqow6 = (Exqow6 & Lxqow6);
assign Lxqow6 = (~(vis_r2_o[29] & Dmqow6));
assign Exqow6 = (~(vis_r6_o[29] & Kmqow6));
assign Qwqow6 = (Sxqow6 & Zxqow6);
assign Zxqow6 = (~(vis_r5_o[29] & Fnqow6));
assign Sxqow6 = (~(vis_r4_o[29] & Mnqow6));
assign Cwqow6 = (Gyqow6 & Nyqow6);
assign Nyqow6 = (Uyqow6 & Bzqow6);
assign Bzqow6 = (~(vis_r1_o[29] & Voqow6));
assign Uyqow6 = (~(vis_r0_o[29] & Cpqow6));
assign Gyqow6 = (Izqow6 & Pzqow6);
assign Pzqow6 = (~(vis_r3_o[29] & Xpqow6));
assign Izqow6 = (~(vis_r7_o[29] & Eqqow6));
assign Lqqow6 = (Wzqow6 & D0row6);
assign D0row6 = (~(K0row6 & Sz8ju6));
assign Wzqow6 = (~(M94iu6 & R0nhu6));
assign M94iu6 = (Shhpw6[29] & Iqzhu6);
assign Jbqow6 = (~(HWDATA[30] | HWDATA[31]));
assign Vaqow6 = (R0row6 & Y0row6);
assign Y0row6 = (~(HWDATA[27] | HWDATA[28]));
assign R0row6 = (~(HWDATA[18] | HWDATA[25]));
assign Haqow6 = (F1row6 & M1row6);
assign M1row6 = (T1row6 & A2row6);
assign A2row6 = (HWDATA[24] & HWDATA[26]);
assign T1row6 = (HWDATA[22] & HWDATA[23]);
assign F1row6 = (H2row6 & O2row6);
assign O2row6 = (HWDATA[20] & HWDATA[21]);
assign H2row6 = (HWDATA[17] & HWDATA[19]);
assign Raohu6 = (Eh6iu6 ? Qnghu6 : V2row6);
assign Eh6iu6 = (!HREADY);
assign V2row6 = (C3row6 & J3row6);
assign J3row6 = (Q3row6 & Udpiu6);
assign Udpiu6 = (!Pzwiu6);
assign Q3row6 = (~(Stdhu6 & Gsaiu6));
assign Gsaiu6 = (~(Xe9ow6 & X3row6));
assign X3row6 = (~(E4row6 & Y2oiu6));
assign E4row6 = (Iugiu6 | P8oiu6);
assign P8oiu6 = (~(Et0ju6 | Xe8iu6));
assign Et0ju6 = (Nlaiu6 | K9aiu6);
assign C3row6 = (U6piu6 & Usaiu6);
assign Usaiu6 = (~(Qa5iu6 | L4row6));
assign L4row6 = (Fsdhu6 & Ja5iu6);
assign Ja5iu6 = (S4row6 & Sf7ju6);
assign Sf7ju6 = (Z4row6 & F23ju6);
assign Z4row6 = (~(As0iu6 | H4ghu6));
assign S4row6 = (Pt2ju6 & Cyfpw6[3]);
assign Qa5iu6 = (Su8ow6 & Xe9ow6);
assign Xe9ow6 = (~(Iepiu6 & Cyfpw6[5]));
assign Su8ow6 = (~(Vo3ju6 & G5row6));
assign G5row6 = (~(N5row6 & U5row6));
assign U5row6 = (~(B6row6 & X97ow6));
assign B6row6 = (Qe8iu6 & Tfjiu6);
assign N5row6 = (~(N4kiu6 & Hs0iu6));
assign N4kiu6 = (I6row6 & Frziu6);
assign I6row6 = (~(Ae0iu6 | C0ehu6));
assign U6piu6 = (P6row6 & Zl1ju6);
assign Zl1ju6 = (~(Emfiu6 & W6row6));
assign W6row6 = (~(D7row6 & Te6iu6));
assign Te6iu6 = (!Ahghu6);
assign D7row6 = (X7gow6 | M2biu6);
assign X7gow6 = (!Righu6);
assign P6row6 = (K7row6 | Sl1ju6);
assign Sl1ju6 = (~(R7row6 & Knbow6));
assign Knbow6 = (Emfiu6 & Y7row6);
assign Y7row6 = (!M2biu6);
assign M2biu6 = (F8row6 & M8row6);
assign Emfiu6 = (~(T8row6 & A9row6));
assign T8row6 = (H9row6 & M8row6);
assign R7row6 = (O9row6 & V0fow6);
assign V0fow6 = (V9row6 | Carow6);
assign V9row6 = (~(Jarow6 & Qarow6));
assign Jarow6 = (~(Ikghu6 & Jhqiu6));
assign O9row6 = (~(Xarow6 & Ebrow6));
assign Ebrow6 = (Lbrow6 | Sbrow6);
assign Xarow6 = (Zbrow6 & Gcrow6);
assign Zbrow6 = (~(Ncrow6 & Ucrow6));
assign Ucrow6 = (Bdrow6 & Idrow6);
assign Bdrow6 = (Okgow6 | Pdrow6);
assign Pdrow6 = (!L1gpw6[0]);
assign Okgow6 = (A8low6 | Wdrow6);
assign Ncrow6 = (~(Derow6 | Kerow6));
assign Kerow6 = (Sbrow6 & Lbrow6);
assign Lbrow6 = (A8low6 ? Yerow6 : Rerow6);
assign Derow6 = (A8low6 ? Mfrow6 : Ffrow6);
assign A8low6 = (~(Tfrow6 & Agrow6));
assign Agrow6 = (~(Carow6 & Hgrow6));
assign Hgrow6 = (~(Ogrow6 & Vgrow6));
assign Vgrow6 = (~(Chrow6 & Jhrow6));
assign Jhrow6 = (Qarow6 ? L1gpw6[0] : B3gpw6[0]);
assign Chrow6 = (~(Mfrow6 | Qhrow6));
assign Qhrow6 = (~(Rerow6 | Xhrow6));
assign Ogrow6 = (~(Xhrow6 & Rerow6));
assign Rerow6 = (Wdrow6 ? B3gpw6[1] : L1gpw6[1]);
assign Xhrow6 = (!Yerow6);
assign Yerow6 = (O8low6 ? Eirow6 : H8gpw6[1]);
assign Carow6 = (~(O8low6 & Lirow6));
assign Lirow6 = (~(Sirow6 & Jhqiu6));
assign Tfrow6 = (Ikghu6 | Wdrow6);
assign Wdrow6 = (!Qarow6);
assign Mfrow6 = (O8low6 ? Zirow6 : H8gpw6[0]);
assign O8low6 = (~(Gjrow6 & Yyghu6));
assign Gjrow6 = (Njrow6 & Jhqiu6);
assign Njrow6 = (~(Sirow6 & Ujrow6));
assign Ujrow6 = (~(Bkrow6 & Ikrow6));
assign Ikrow6 = (Pkrow6 | Zirow6);
assign Pkrow6 = (~(H8gpw6[0] & Wkrow6));
assign Wkrow6 = (Dlrow6 | H8gpw6[1]);
assign Bkrow6 = (~(H8gpw6[1] & Dlrow6));
assign Dlrow6 = (!Eirow6);
assign Eirow6 = (E2fow6 ? Rlrow6 : Klrow6);
assign Klrow6 = (!Ylrow6);
assign Sirow6 = (~(Fmrow6 & Mmrow6));
assign Mmrow6 = (~(E2fow6 | H7fow6));
assign E2fow6 = (!Meeow6);
assign Fmrow6 = (C8fow6 & Tmrow6);
assign Zirow6 = (Meeow6 ? Hnrow6 : Anrow6);
assign Meeow6 = (~(Onrow6 & Vnrow6));
assign Vnrow6 = (~(Corow6 & Jorow6));
assign Jorow6 = (Ylrow6 | Rlrow6);
assign Corow6 = (Qorow6 & Xorow6);
assign Xorow6 = (~(Eprow6 & C8fow6));
assign Eprow6 = (Tmrow6 & Lprow6);
assign Qorow6 = (~(Sprow6 & Zprow6));
assign Zprow6 = (~(Rlrow6 & Ylrow6));
assign Ylrow6 = (H7fow6 ? Nqrow6 : Gqrow6);
assign Nqrow6 = (!Uqrow6);
assign Rlrow6 = (B4fow6 ? Irrow6 : Brrow6);
assign Brrow6 = (!Prrow6);
assign Sprow6 = (Hnrow6 | Wrrow6);
assign Wrrow6 = (!Anrow6);
assign Onrow6 = (Dsrow6 | B4fow6);
assign Hnrow6 = (Ksrow6 | Rsrow6);
assign Rsrow6 = (~(F6fow6 | Ysrow6));
assign F6fow6 = (Lprow6 | Ftrow6);
assign Ksrow6 = (H7fow6 ? Ttrow6 : Mtrow6);
assign H7fow6 = (!Lprow6);
assign Lprow6 = (~(Aurow6 & Hurow6));
assign Hurow6 = (~(Ourow6 & Vurow6));
assign Vurow6 = (~(Cvrow6 & Jvrow6));
assign Jvrow6 = (~(Uqrow6 & Gqrow6));
assign Cvrow6 = (~(Qvrow6 & Xvrow6));
assign Xvrow6 = (O7fow6 ? Lwrow6 : Ewrow6);
assign Qvrow6 = (~(Mtrow6 | Swrow6));
assign Swrow6 = (~(Gqrow6 | Uqrow6));
assign Uqrow6 = (Ftrow6 ? Gxrow6 : Zwrow6);
assign Gqrow6 = (Hdgow6 ? Uxrow6 : Nxrow6);
assign Ourow6 = (~(C8fow6 & Tmrow6));
assign C8fow6 = (Q8fow6 & Jegow6);
assign Aurow6 = (~(Byrow6 & Iyrow6));
assign Byrow6 = (~(Pyrow6 | Ftrow6));
assign Ttrow6 = (Ftrow6 & Ewrow6);
assign Ftrow6 = (!O7fow6);
assign O7fow6 = (~(Wyrow6 & Dzrow6));
assign Dzrow6 = (~(Kzrow6 & Rzrow6));
assign Rzrow6 = (Yzrow6 | Gxrow6);
assign Kzrow6 = (F0sow6 & M0sow6);
assign M0sow6 = (~(Iyrow6 & T0sow6));
assign T0sow6 = (!Pyrow6);
assign Iyrow6 = (~(M6fow6 | A1sow6));
assign F0sow6 = (~(H1sow6 & O1sow6));
assign O1sow6 = (~(Gxrow6 & Yzrow6));
assign Yzrow6 = (!Zwrow6);
assign Zwrow6 = (M6fow6 ? C2sow6 : V1sow6);
assign Gxrow6 = (X2sow6 ? Q2sow6 : J2sow6);
assign H1sow6 = (~(Ysrow6 & Ewrow6));
assign Ewrow6 = (V7fow6 ? L3sow6 : E3sow6);
assign V7fow6 = (!X2sow6);
assign Ysrow6 = (!Lwrow6);
assign Lwrow6 = (M6fow6 ? Z3sow6 : S3sow6);
assign M6fow6 = (G4sow6 & N4sow6);
assign N4sow6 = (~(U4sow6 & B5sow6));
assign B5sow6 = (~(I5sow6 & P5sow6));
assign P5sow6 = (W5sow6 | D6sow6);
assign D6sow6 = (Wagow6 ? R4gpw6[46] : R4gpw6[44]);
assign W5sow6 = (~(Z3sow6 & K6sow6));
assign K6sow6 = (~(V1sow6 & R6sow6));
assign I5sow6 = (R6sow6 | V1sow6);
assign V1sow6 = (Wagow6 ? R4gpw6[47] : R4gpw6[45]);
assign Wagow6 = (!A1sow6);
assign R6sow6 = (!C2sow6);
assign C2sow6 = (Dbgow6 ? R4gpw6[43] : R4gpw6[41]);
assign U4sow6 = (Pyrow6 | A1sow6);
assign G4sow6 = (~(Dbgow6 & Y6sow6));
assign Y6sow6 = (~(Vbgpw6[21] & Odgpw6[21]));
assign Z3sow6 = (F7sow6 ? R4gpw6[40] : R4gpw6[42]);
assign F7sow6 = (!Dbgow6);
assign Dbgow6 = (~(M7sow6 & Vbgpw6[20]));
assign M7sow6 = (Odgpw6[20] & T7sow6);
assign T7sow6 = (~(A8sow6 & Vbgpw6[21]));
assign A8sow6 = (Odgpw6[21] & H8sow6);
assign H8sow6 = (~(O8sow6 & V8sow6));
assign V8sow6 = (~(C9sow6 & R4gpw6[40]));
assign C9sow6 = (~(J9sow6 | R4gpw6[42]));
assign J9sow6 = (~(Q9sow6 | R4gpw6[41]));
assign O8sow6 = (~(R4gpw6[41] & Q9sow6));
assign S3sow6 = (A1sow6 ? R4gpw6[44] : R4gpw6[46]);
assign A1sow6 = (X9sow6 & Vbgpw6[22]);
assign X9sow6 = (Odgpw6[22] & Easow6);
assign Easow6 = (~(Lasow6 & Pyrow6));
assign Pyrow6 = (Vbgpw6[23] & Odgpw6[23]);
assign Lasow6 = (Sasow6 & Zasow6);
assign Zasow6 = (~(Gbsow6 & Nbsow6));
assign Nbsow6 = (Ubsow6 | R4gpw6[47]);
assign Gbsow6 = (~(R4gpw6[44] & Bcsow6));
assign Sasow6 = (~(R4gpw6[47] & Ubsow6));
assign Wyrow6 = (~(Icsow6 & Pcsow6));
assign Icsow6 = (X2sow6 & Kbgow6);
assign X2sow6 = (~(Wcsow6 & Ddsow6));
assign Ddsow6 = (~(Kdsow6 & Rdsow6));
assign Rdsow6 = (~(Ydsow6 & Fesow6));
assign Fesow6 = (~(Mesow6 & L3sow6));
assign L3sow6 = (Rbgow6 ? R4gpw6[34] : R4gpw6[32]);
assign Mesow6 = (~(E3sow6 | Tesow6));
assign Tesow6 = (~(Afsow6 | J2sow6));
assign E3sow6 = (Kbgow6 ? R4gpw6[38] : R4gpw6[36]);
assign Ydsow6 = (~(J2sow6 & Afsow6));
assign Afsow6 = (!Q2sow6);
assign Q2sow6 = (Kbgow6 ? R4gpw6[39] : R4gpw6[37]);
assign J2sow6 = (Rbgow6 ? R4gpw6[35] : R4gpw6[33]);
assign Kdsow6 = (~(Pcsow6 & Kbgow6));
assign Kbgow6 = (~(Hfsow6 & Vbgpw6[18]));
assign Hfsow6 = (Odgpw6[18] & Ofsow6);
assign Ofsow6 = (Vfsow6 | Pcsow6);
assign Vfsow6 = (~(Cgsow6 & Jgsow6));
assign Jgsow6 = (~(Qgsow6 & Xgsow6));
assign Xgsow6 = (Ehsow6 | R4gpw6[39]);
assign Qgsow6 = (~(R4gpw6[36] & Lhsow6));
assign Cgsow6 = (~(R4gpw6[39] & Ehsow6));
assign Pcsow6 = (~(Vbgpw6[19] & Odgpw6[19]));
assign Wcsow6 = (~(Rbgow6 & Shsow6));
assign Shsow6 = (~(Vbgpw6[17] & Odgpw6[17]));
assign Rbgow6 = (~(Zhsow6 & Vbgpw6[16]));
assign Zhsow6 = (Odgpw6[16] & Gisow6);
assign Gisow6 = (~(Nisow6 & Uisow6));
assign Uisow6 = (Bjsow6 & Ijsow6);
assign Ijsow6 = (~(Pjsow6 & Wjsow6));
assign Wjsow6 = (~(R4gpw6[33] & Dksow6));
assign Pjsow6 = (~(R4gpw6[32] & Kksow6));
assign Kksow6 = (!R4gpw6[34]);
assign Bjsow6 = (Dksow6 | R4gpw6[33]);
assign Nisow6 = (Vbgpw6[17] & Odgpw6[17]);
assign Mtrow6 = (Hdgow6 ? Yksow6 : Rksow6);
assign Hdgow6 = (!Q8fow6);
assign Q8fow6 = (~(Flsow6 & Mlsow6));
assign Mlsow6 = (Tlsow6 | Amsow6);
assign Tlsow6 = (X8fow6 | Vdgow6);
assign Flsow6 = (~(Hmsow6 & Omsow6));
assign Omsow6 = (~(Vmsow6 & Cnsow6));
assign Cnsow6 = (~(Jnsow6 & Qnsow6));
assign Qnsow6 = (Xnsow6 & Eosow6);
assign Xnsow6 = (Nxrow6 | Losow6);
assign Jnsow6 = (Yksow6 & Sosow6);
assign Vmsow6 = (~(Losow6 & Nxrow6));
assign Nxrow6 = (Jegow6 ? Gpsow6 : Zosow6);
assign Zosow6 = (!Npsow6);
assign Losow6 = (!Uxrow6);
assign Uxrow6 = (X8fow6 ? Bqsow6 : Upsow6);
assign X8fow6 = (!Cegow6);
assign Hmsow6 = (~(Tmrow6 & Jegow6));
assign Yksow6 = (Cegow6 ? Pqsow6 : Iqsow6);
assign Cegow6 = (~(Wqsow6 & Drsow6));
assign Drsow6 = (~(Krsow6 & Rrsow6));
assign Rrsow6 = (~(Yrsow6 & Fssow6));
assign Fssow6 = (~(Mssow6 & Iqsow6));
assign Mssow6 = (~(Pqsow6 | Tssow6));
assign Tssow6 = (~(Atsow6 | Upsow6));
assign Yrsow6 = (~(Upsow6 & Atsow6));
assign Atsow6 = (!Bqsow6);
assign Bqsow6 = (Odgow6 ? Otsow6 : Htsow6);
assign Upsow6 = (Jusow6 ? Cusow6 : Vtsow6);
assign Krsow6 = (Amsow6 | Vdgow6);
assign Wqsow6 = (Odgow6 | Qusow6);
assign Pqsow6 = (Jusow6 ? R4gpw6[54] : R4gpw6[52]);
assign Jusow6 = (!Vdgow6);
assign Vdgow6 = (Xusow6 & Vbgpw6[26]);
assign Xusow6 = (Odgpw6[26] & Evsow6);
assign Evsow6 = (~(Lvsow6 & Amsow6));
assign Amsow6 = (Vbgpw6[27] & Odgpw6[27]);
assign Lvsow6 = (Svsow6 & Zvsow6);
assign Zvsow6 = (~(Gwsow6 & Nwsow6));
assign Nwsow6 = (Vtsow6 | R4gpw6[55]);
assign Gwsow6 = (Uwsow6 | R4gpw6[54]);
assign Svsow6 = (Cusow6 | R4gpw6[53]);
assign Iqsow6 = (Odgow6 ? R4gpw6[48] : R4gpw6[50]);
assign Odgow6 = (Bxsow6 & Vbgpw6[24]);
assign Bxsow6 = (Odgpw6[24] & Ixsow6);
assign Ixsow6 = (~(Qusow6 & Pxsow6));
assign Pxsow6 = (Wxsow6 & Dysow6);
assign Dysow6 = (~(Kysow6 & Rysow6));
assign Rysow6 = (Otsow6 | R4gpw6[51]);
assign Kysow6 = (Yysow6 | R4gpw6[50]);
assign Wxsow6 = (Htsow6 | R4gpw6[49]);
assign Qusow6 = (Vbgpw6[25] & Odgpw6[25]);
assign Rksow6 = (~(Eosow6 & Sosow6));
assign Sosow6 = (~(Fzsow6 & Jegow6));
assign Eosow6 = (~(Mzsow6 & Tzsow6));
assign Mzsow6 = (!Jegow6);
assign Jegow6 = (~(A0tow6 & H0tow6));
assign H0tow6 = (Tmrow6 | O0tow6);
assign O0tow6 = (V0tow6 & C1tow6);
assign C1tow6 = (~(J1tow6 & Tzsow6));
assign Tzsow6 = (Q1tow6 ? R4gpw6[58] : R4gpw6[56]);
assign J1tow6 = (~(Fzsow6 | X1tow6));
assign X1tow6 = (~(Npsow6 | Gpsow6));
assign Fzsow6 = (Mcgow6 ? R4gpw6[62] : R4gpw6[60]);
assign V0tow6 = (~(Gpsow6 & Npsow6));
assign Npsow6 = (Qegow6 ? R4gpw6[57] : R4gpw6[59]);
assign Qegow6 = (!Q1tow6);
assign Gpsow6 = (Mcgow6 ? L2tow6 : E2tow6);
assign Tmrow6 = (Mcgow6 & S2tow6);
assign S2tow6 = (~(Vbgpw6[31] & Odgpw6[31]));
assign Mcgow6 = (~(Z2tow6 & Vbgpw6[30]));
assign Z2tow6 = (Odgpw6[30] & G3tow6);
assign G3tow6 = (~(N3tow6 & U3tow6));
assign U3tow6 = (B4tow6 & I4tow6);
assign I4tow6 = (~(P4tow6 & W4tow6));
assign W4tow6 = (E2tow6 | R4gpw6[63]);
assign P4tow6 = (~(R4gpw6[60] & D5tow6));
assign D5tow6 = (!R4gpw6[62]);
assign B4tow6 = (L2tow6 | R4gpw6[61]);
assign L2tow6 = (!R4gpw6[63]);
assign N3tow6 = (Vbgpw6[31] & Odgpw6[31]);
assign A0tow6 = (~(Q1tow6 & K5tow6));
assign K5tow6 = (~(Vbgpw6[29] & Odgpw6[29]));
assign Q1tow6 = (~(R5tow6 & Vbgpw6[28]));
assign R5tow6 = (Odgpw6[28] & Y5tow6);
assign Y5tow6 = (~(F6tow6 & Vbgpw6[29]));
assign F6tow6 = (Odgpw6[29] & M6tow6);
assign M6tow6 = (~(T6tow6 & A7tow6));
assign A7tow6 = (~(H7tow6 & R4gpw6[56]));
assign H7tow6 = (~(O7tow6 | R4gpw6[58]));
assign O7tow6 = (~(V7tow6 | R4gpw6[57]));
assign T6tow6 = (~(R4gpw6[57] & V7tow6));
assign Anrow6 = (~(C8tow6 & J8tow6));
assign J8tow6 = (~(Z2fow6 & Q8tow6));
assign Q8tow6 = (~(X8tow6 & E9tow6));
assign Z2fow6 = (B4fow6 & I4fow6);
assign C8tow6 = (B4fow6 ? S9tow6 : L9tow6);
assign B4fow6 = (!Sfgow6);
assign Sfgow6 = (~(Z9tow6 & Gatow6));
assign Gatow6 = (~(Dsrow6 & Natow6));
assign Natow6 = (~(Uatow6 & Bbtow6));
assign Bbtow6 = (~(Ibtow6 & Pbtow6));
assign Pbtow6 = (Wbtow6 & Dctow6);
assign Wbtow6 = (Prrow6 | Irrow6);
assign Ibtow6 = (~(Kctow6 | Rctow6));
assign Rctow6 = (Nggow6 & Yctow6);
assign Kctow6 = (Yigow6 ? Mdtow6 : Fdtow6);
assign Uatow6 = (~(Irrow6 & Prrow6));
assign Prrow6 = (Nggow6 ? Aetow6 : Tdtow6);
assign Irrow6 = (Yigow6 ? Oetow6 : Hetow6);
assign Dsrow6 = (~(Vetow6 & Cftow6));
assign Vetow6 = (~(Jftow6 | Nggow6));
assign Z9tow6 = (~(Qftow6 & Xftow6));
assign Qftow6 = (~(Egtow6 | Yigow6));
assign Yigow6 = (!I4fow6);
assign S9tow6 = (I4fow6 | Mdtow6);
assign Mdtow6 = (!Lgtow6);
assign I4fow6 = (~(Sgtow6 & Zgtow6));
assign Zgtow6 = (Ghtow6 | Nhtow6);
assign Ghtow6 = (P4fow6 | Mjgow6);
assign Sgtow6 = (~(Uhtow6 & Bitow6));
assign Bitow6 = (~(Xftow6 & Iitow6));
assign Iitow6 = (!Egtow6);
assign Xftow6 = (~(Pitow6 | Hkgow6));
assign Uhtow6 = (~(Witow6 & Djtow6));
assign Djtow6 = (~(Kjtow6 & Fdtow6));
assign Fdtow6 = (X8tow6 & E9tow6);
assign E9tow6 = (~(Pitow6 & Rjtow6));
assign X8tow6 = (~(Yjtow6 & G3fow6));
assign Kjtow6 = (Lgtow6 & Fktow6);
assign Fktow6 = (Mktow6 | Oetow6);
assign Lgtow6 = (P4fow6 ? Altow6 : Tktow6);
assign P4fow6 = (!Tjgow6);
assign Altow6 = (Fjgow6 ? R4gpw6[0] : R4gpw6[2]);
assign Witow6 = (~(Oetow6 & Mktow6));
assign Mktow6 = (!Hetow6);
assign Hetow6 = (Pitow6 ? Oltow6 : Hltow6);
assign Pitow6 = (!G3fow6);
assign G3fow6 = (~(Vltow6 & Cmtow6));
assign Cmtow6 = (~(Jmtow6 & Qmtow6));
assign Qmtow6 = (~(Xmtow6 & Entow6));
assign Entow6 = (~(Lntow6 & Rjtow6));
assign Rjtow6 = (Akgow6 ? R4gpw6[8] : R4gpw6[10]);
assign Lntow6 = (~(Yjtow6 | Sntow6));
assign Sntow6 = (~(Zntow6 | Oltow6));
assign Yjtow6 = (Hkgow6 ? R4gpw6[12] : R4gpw6[14]);
assign Xmtow6 = (~(Oltow6 & Zntow6));
assign Jmtow6 = (Egtow6 | Hkgow6);
assign Vltow6 = (~(Gotow6 & Notow6));
assign Notow6 = (~(Vbgpw6[5] & Odgpw6[5]));
assign Oltow6 = (Akgow6 ? R4gpw6[9] : R4gpw6[11]);
assign Akgow6 = (!Gotow6);
assign Gotow6 = (~(Uotow6 & Vbgpw6[4]));
assign Uotow6 = (Odgpw6[4] & Bptow6);
assign Bptow6 = (~(Iptow6 & Vbgpw6[5]));
assign Iptow6 = (Odgpw6[5] & Pptow6);
assign Pptow6 = (~(Wptow6 & Dqtow6));
assign Dqtow6 = (~(Kqtow6 & R4gpw6[8]));
assign Kqtow6 = (~(Rqtow6 | R4gpw6[10]));
assign Rqtow6 = (~(Yqtow6 | R4gpw6[9]));
assign Wptow6 = (~(R4gpw6[9] & Yqtow6));
assign Hltow6 = (!Zntow6);
assign Zntow6 = (Hkgow6 ? Mrtow6 : Frtow6);
assign Hkgow6 = (Trtow6 & Vbgpw6[6]);
assign Trtow6 = (Odgpw6[6] & Astow6);
assign Astow6 = (~(Hstow6 & Egtow6));
assign Egtow6 = (Vbgpw6[7] & Odgpw6[7]);
assign Hstow6 = (Ostow6 & Vstow6);
assign Vstow6 = (~(Cttow6 & Jttow6));
assign Jttow6 = (Mrtow6 | R4gpw6[15]);
assign Cttow6 = (~(R4gpw6[12] & Qttow6));
assign Ostow6 = (Frtow6 | R4gpw6[13]);
assign Oetow6 = (Tjgow6 ? Eutow6 : Xttow6);
assign Tjgow6 = (~(Lutow6 & Sutow6));
assign Sutow6 = (~(Zutow6 & Gvtow6));
assign Gvtow6 = (~(Nvtow6 & Uvtow6));
assign Uvtow6 = (~(Bwtow6 & Iwtow6));
assign Iwtow6 = (Pwtow6 ? R4gpw6[2] : R4gpw6[0]);
assign Bwtow6 = (~(Tktow6 | Wwtow6));
assign Wwtow6 = (~(Dxtow6 | Xttow6));
assign Tktow6 = (Kxtow6 ? R4gpw6[6] : R4gpw6[4]);
assign Kxtow6 = (!Mjgow6);
assign Nvtow6 = (~(Xttow6 & Dxtow6));
assign Zutow6 = (Nhtow6 | Mjgow6);
assign Lutow6 = (~(Pwtow6 & Rxtow6));
assign Rxtow6 = (~(Vbgpw6[1] & Odgpw6[1]));
assign Eutow6 = (!Dxtow6);
assign Dxtow6 = (Mjgow6 ? Fytow6 : Yxtow6);
assign Mjgow6 = (Mytow6 & Vbgpw6[2]);
assign Mytow6 = (Odgpw6[2] & Tytow6);
assign Tytow6 = (~(Aztow6 & Nhtow6));
assign Nhtow6 = (Vbgpw6[3] & Odgpw6[3]);
assign Aztow6 = (Hztow6 & Oztow6);
assign Oztow6 = (~(Vztow6 & C0uow6));
assign C0uow6 = (Fytow6 | R4gpw6[7]);
assign Vztow6 = (J0uow6 | R4gpw6[6]);
assign Hztow6 = (Yxtow6 | R4gpw6[5]);
assign Xttow6 = (Fjgow6 ? R4gpw6[1] : R4gpw6[3]);
assign Fjgow6 = (!Pwtow6);
assign Pwtow6 = (~(Q0uow6 & Vbgpw6[0]));
assign Q0uow6 = (Odgpw6[0] & X0uow6);
assign X0uow6 = (~(E1uow6 & L1uow6));
assign L1uow6 = (S1uow6 & Z1uow6);
assign Z1uow6 = (~(G2uow6 & N2uow6));
assign N2uow6 = (U2uow6 | R4gpw6[3]);
assign G2uow6 = (B3uow6 | R4gpw6[2]);
assign S1uow6 = (~(R4gpw6[3] & U2uow6));
assign E1uow6 = (Vbgpw6[1] & Odgpw6[1]);
assign L9tow6 = (I3uow6 & Dctow6);
assign Dctow6 = (~(K5fow6 & P3uow6));
assign P3uow6 = (~(W3uow6 & D4uow6));
assign I3uow6 = (~(Nggow6 & Yctow6));
assign Nggow6 = (!K5fow6);
assign K5fow6 = (~(K4uow6 & R4uow6));
assign R4uow6 = (Y4uow6 | F5uow6);
assign Y4uow6 = (W4fow6 | Bhgow6);
assign K4uow6 = (~(M5uow6 & T5uow6));
assign T5uow6 = (~(Cftow6 & A6uow6));
assign A6uow6 = (!Jftow6);
assign Cftow6 = (~(D5fow6 | Whgow6));
assign M5uow6 = (~(H6uow6 & O6uow6));
assign O6uow6 = (~(V6uow6 & C7uow6));
assign C7uow6 = (J7uow6 & D4uow6);
assign D4uow6 = (~(D5fow6 & Q7uow6));
assign D5fow6 = (!Digow6);
assign J7uow6 = (Tdtow6 | X7uow6);
assign V6uow6 = (Yctow6 & W3uow6);
assign W3uow6 = (~(E8uow6 & Digow6));
assign Yctow6 = (W4fow6 ? S8uow6 : L8uow6);
assign S8uow6 = (Uggow6 ? R4gpw6[16] : R4gpw6[18]);
assign H6uow6 = (~(X7uow6 & Tdtow6));
assign Tdtow6 = (Digow6 ? G9uow6 : Z8uow6);
assign Digow6 = (~(N9uow6 & U9uow6));
assign U9uow6 = (~(Bauow6 & Iauow6));
assign Iauow6 = (~(Pauow6 & Wauow6));
assign Wauow6 = (~(Dbuow6 & Q7uow6));
assign Q7uow6 = (Phgow6 ? R4gpw6[24] : R4gpw6[26]);
assign Dbuow6 = (~(E8uow6 | Kbuow6));
assign Kbuow6 = (~(G9uow6 | Rbuow6));
assign E8uow6 = (Whgow6 ? R4gpw6[28] : R4gpw6[30]);
assign Pauow6 = (~(Rbuow6 & G9uow6));
assign Bauow6 = (Jftow6 | Whgow6);
assign N9uow6 = (~(Ybuow6 & Fcuow6));
assign Fcuow6 = (~(Vbgpw6[13] & Odgpw6[13]));
assign G9uow6 = (Whgow6 ? Tcuow6 : Mcuow6);
assign Whgow6 = (Aduow6 & Vbgpw6[14]);
assign Aduow6 = (Odgpw6[14] & Hduow6);
assign Hduow6 = (~(Oduow6 & Jftow6));
assign Jftow6 = (Vbgpw6[15] & Odgpw6[15]);
assign Oduow6 = (Vduow6 & Ceuow6);
assign Ceuow6 = (~(Jeuow6 & Qeuow6));
assign Qeuow6 = (Tcuow6 | R4gpw6[31]);
assign Jeuow6 = (~(R4gpw6[28] & Xeuow6));
assign Xeuow6 = (!R4gpw6[30]);
assign Vduow6 = (Mcuow6 | R4gpw6[29]);
assign Tcuow6 = (!R4gpw6[29]);
assign Z8uow6 = (!Rbuow6);
assign Rbuow6 = (Phgow6 ? R4gpw6[25] : R4gpw6[27]);
assign Phgow6 = (!Ybuow6);
assign Ybuow6 = (~(Efuow6 & Vbgpw6[12]));
assign Efuow6 = (Odgpw6[12] & Lfuow6);
assign Lfuow6 = (~(Sfuow6 & Vbgpw6[13]));
assign Sfuow6 = (Odgpw6[13] & Zfuow6);
assign Zfuow6 = (~(Gguow6 & Nguow6));
assign Nguow6 = (~(Uguow6 & R4gpw6[24]));
assign Uguow6 = (~(Bhuow6 | R4gpw6[26]));
assign Bhuow6 = (~(Ihuow6 | R4gpw6[25]));
assign Gguow6 = (~(R4gpw6[25] & Ihuow6));
assign X7uow6 = (!Aetow6);
assign Aetow6 = (W4fow6 ? Whuow6 : Phuow6);
assign W4fow6 = (!Ihgow6);
assign Ihgow6 = (~(Diuow6 & Kiuow6));
assign Kiuow6 = (~(Riuow6 & Yiuow6));
assign Yiuow6 = (~(Fjuow6 & Mjuow6));
assign Mjuow6 = (~(Tjuow6 & Akuow6));
assign Akuow6 = (Hkuow6 ? R4gpw6[18] : R4gpw6[16]);
assign Tjuow6 = (~(L8uow6 | Okuow6));
assign Okuow6 = (~(Vkuow6 | Phuow6));
assign L8uow6 = (Cluow6 ? R4gpw6[22] : R4gpw6[20]);
assign Fjuow6 = (~(Phuow6 & Vkuow6));
assign Vkuow6 = (!Whuow6);
assign Riuow6 = (F5uow6 | Bhgow6);
assign Diuow6 = (~(Hkuow6 & Jluow6));
assign Jluow6 = (~(Vbgpw6[9] & Odgpw6[9]));
assign Whuow6 = (Uggow6 ? Xluow6 : Qluow6);
assign Uggow6 = (!Hkuow6);
assign Hkuow6 = (~(Emuow6 & Vbgpw6[8]));
assign Emuow6 = (Odgpw6[8] & Lmuow6);
assign Lmuow6 = (~(Smuow6 & Zmuow6));
assign Zmuow6 = (Gnuow6 & Nnuow6);
assign Nnuow6 = (~(Unuow6 & Bouow6));
assign Bouow6 = (Xluow6 | R4gpw6[19]);
assign Unuow6 = (Iouow6 | R4gpw6[18]);
assign Gnuow6 = (Qluow6 | R4gpw6[17]);
assign Smuow6 = (Vbgpw6[9] & Odgpw6[9]);
assign Phuow6 = (Cluow6 ? Wouow6 : Pouow6);
assign Cluow6 = (!Bhgow6);
assign Bhgow6 = (Dpuow6 & Vbgpw6[10]);
assign Dpuow6 = (Odgpw6[10] & Kpuow6);
assign Kpuow6 = (~(Rpuow6 & F5uow6));
assign F5uow6 = (Vbgpw6[11] & Odgpw6[11]);
assign Rpuow6 = (Ypuow6 & Fquow6);
assign Fquow6 = (~(Mquow6 & Tquow6));
assign Tquow6 = (Pouow6 | R4gpw6[23]);
assign Mquow6 = (Aruow6 | R4gpw6[22]);
assign Ypuow6 = (Wouow6 | R4gpw6[21]);
assign Ffrow6 = (~(Qarow6 | Xglow6));
assign Qarow6 = (~(Zlghu6 & Hruow6));
assign Hruow6 = (~(Oruow6 & Vruow6));
assign Vruow6 = (Csuow6 & Jhqiu6);
assign Jhqiu6 = (~(P9hhu6 & Jehhu6));
assign Csuow6 = (~(Jsuow6 & Qsuow6));
assign Qsuow6 = (F4oow6 | L1gpw6[1]);
assign Jsuow6 = (Xglow6 | L1gpw6[0]);
assign Oruow6 = (Ikghu6 & Xsuow6);
assign Xsuow6 = (~(L1gpw6[1] & F4oow6));
assign F4oow6 = (!B3gpw6[1]);
assign K7row6 = (Cz8iu6 ? vis_primask_o : Oy8iu6);
assign Cz8iu6 = (Etuow6 & Ltuow6);
assign Ltuow6 = (~(Stuow6 & Ztuow6));
assign Ztuow6 = (Cyfpw6[4] & Gmniu6);
assign Gmniu6 = (~(Guuow6 & Nuuow6));
assign Nuuow6 = (Uuuow6 & Bvuow6);
assign Bvuow6 = (Ivuow6 | Yoniu6);
assign Yoniu6 = (Pvuow6 & Wvuow6);
assign Wvuow6 = (~(Dwuow6 & Kwuow6));
assign Dwuow6 = (~(C0ehu6 | H4ghu6));
assign Pvuow6 = (~(Glaiu6 | Rwuow6));
assign Rwuow6 = (Ywuow6 & Fxuow6);
assign Fxuow6 = (~(Nlaiu6 | Hs0iu6));
assign Ywuow6 = (Jf6ju6 & Imaiu6);
assign Uuuow6 = (Mxuow6 | Mpniu6);
assign Mpniu6 = (Txuow6 & Ayuow6);
assign Ayuow6 = (Hyuow6 & Xiaju6);
assign Xiaju6 = (Oyuow6 & W8oiu6);
assign Oyuow6 = (~(Vyuow6 & Ae0iu6));
assign Vyuow6 = (U4kiu6 & Yljiu6);
assign Hyuow6 = (Czuow6 & Jzuow6);
assign Jzuow6 = (Z6oiu6 | E4jiu6);
assign Z6oiu6 = (!Fhaiu6);
assign Czuow6 = (~(Qzuow6 & Cyfpw6[7]));
assign Qzuow6 = (Cyfpw6[1] & Xzuow6);
assign Xzuow6 = (~(E0vow6 & Vwaiu6));
assign E0vow6 = (Y7ghu6 | Cyfpw6[4]);
assign Txuow6 = (L0vow6 & S0vow6);
assign S0vow6 = (Cyfpw6[4] ? G1vow6 : Z0vow6);
assign G1vow6 = (Nlaiu6 | Mr0iu6);
assign Z0vow6 = (Qxaiu6 | Cyfpw6[6]);
assign L0vow6 = (N1vow6 & U1vow6);
assign U1vow6 = (~(Xe8iu6 & B2vow6));
assign B2vow6 = (U4kiu6 | Vboiu6);
assign N1vow6 = (Yn2ju6 | Ii0iu6);
assign Guuow6 = (Utniu6 & I2vow6);
assign I2vow6 = (~(S8fpw6[9] & Wnniu6));
assign Wnniu6 = (~(P2vow6 & W2vow6));
assign W2vow6 = (~(Gz2ju6 | Iugiu6));
assign Gz2ju6 = (~(X5oiu6 | Yn2ju6));
assign Yn2ju6 = (!Pfoiu6);
assign X5oiu6 = (!F9aju6);
assign P2vow6 = (D3vow6 & K3vow6);
assign K3vow6 = (~(R3vow6 & Cyfpw6[4]));
assign R3vow6 = (~(Lkaiu6 | Tr0iu6));
assign D3vow6 = (~(C0ehu6 & Y3vow6));
assign Y3vow6 = (~(F4vow6 & M4vow6));
assign M4vow6 = (G7oiu6 | Hs0iu6);
assign F4vow6 = (T4vow6 & Ekaiu6);
assign Ekaiu6 = (A4oiu6 | Cyfpw6[0]);
assign T4vow6 = (M32ju6 | Tfjiu6);
assign Utniu6 = (~(A5vow6 | Fq8iu6));
assign A5vow6 = (~(Mzlow6 | C0ehu6));
assign Etuow6 = (Vlliu6 & H5vow6);
assign H5vow6 = (~(O5vow6 & Jjoiu6));
assign Jjoiu6 = (B5kiu6 & Qmliu6);
assign B5kiu6 = (!S8fpw6[2]);
assign O5vow6 = (~(Wofiu6 | Qjoiu6));
assign Vlliu6 = (~(V5vow6 & S8fpw6[2]));
assign V5vow6 = (Qmliu6 & Wofiu6);
assign Oy8iu6 = (~(C6vow6 & J6vow6));
assign J6vow6 = (~(Stuow6 & X3fpw6[1]));
assign Stuow6 = (~(M32ju6 | P1bow6));
assign M32ju6 = (!W2aow6);
assign C6vow6 = (~(Qmliu6 & L35ju6));
assign Qmliu6 = (~(Q6vow6 & X6vow6));
assign X6vow6 = (~(E7vow6 & Obbow6));
assign E7vow6 = (~(A4oiu6 | Cyfpw6[6]));
assign A4oiu6 = (!Pugiu6);
assign Q6vow6 = (Kgaiu6 | Ii0iu6);
assign Fmdhu6 = (RSTBYPASS ? PORESETn : Oodhu6);
assign TXEV = (L7vow6 & Iugiu6);
assign Iugiu6 = (S7vow6 & Vo3ju6);
assign S7vow6 = (~(Knaiu6 | Cyfpw6[6]));
assign L7vow6 = (Pt2ju6 & Cyfpw6[4]);
assign SWDO = (Ujyhu6 ? Hknhu6 : Tonhu6);
assign Ujyhu6 = (!Ighpw6[5]);
assign SPECHTRANS = (~(HMASTER & Z7vow6));
assign Z7vow6 = (~(Krzhu6 & Ebxiu6));
assign SLEEPDEEP = (SLEEPING & Ndghu6);
assign HWRITE = (!G8vow6);
assign G8vow6 = (Xg6iu6 ? Sq4iu6 : Ejpiu6);
assign Sq4iu6 = (Iqnhu6 & Iqzhu6);
assign Ejpiu6 = (N8vow6 & U8vow6);
assign U8vow6 = (B9vow6 & I9vow6);
assign I9vow6 = (~(Xzmiu6 & P9vow6));
assign P9vow6 = (W9vow6 | Bi0iu6);
assign Bi0iu6 = (Wp0iu6 & Y7ghu6);
assign W9vow6 = (Kwuow6 & Wp0iu6);
assign Kwuow6 = (~(Qjaiu6 | Xkaow6));
assign B9vow6 = (~(Us2ju6 & Davow6));
assign Davow6 = (Kavow6 | Moaiu6);
assign Moaiu6 = (D6kiu6 & Y2oiu6);
assign Kavow6 = (Ravow6 & Ldoiu6);
assign Ravow6 = (~(P1bow6 | Sbghu6));
assign Us2ju6 = (Cyfpw6[7] & Gwyiu6);
assign N8vow6 = (Lv7ow6 & Yavow6);
assign Lv7ow6 = (Fbvow6 & Oe8ow6);
assign Fbvow6 = (~(Mbvow6 & Ldoiu6));
assign Mbvow6 = (Qe8iu6 & H4ghu6);
assign HWDATA[9] = (~(Tbvow6 & Acvow6));
assign Tbvow6 = (Hcvow6 & Ocvow6);
assign Ocvow6 = (~(Ym4iu6 & R0nhu6));
assign Ym4iu6 = (Shhpw6[9] & Iqzhu6);
assign Hcvow6 = (Vcvow6 | I28ju6);
assign HWDATA[8] = (~(Cdvow6 & Jdvow6));
assign Cdvow6 = (Qdvow6 & Xdvow6);
assign Xdvow6 = (~(Pl4iu6 & R0nhu6));
assign Pl4iu6 = (Shhpw6[8] & Iqzhu6);
assign Qdvow6 = (Vcvow6 | Cz7ju6);
assign HWDATA[7] = (~(Eevow6 & Levow6));
assign Levow6 = (~(Gk4iu6 & R0nhu6));
assign Gk4iu6 = (Shhpw6[7] & Iqzhu6);
assign Eevow6 = (~(Sevow6 & Uo6ju6));
assign HWDATA[6] = (~(Zevow6 & Gfvow6));
assign Gfvow6 = (~(Xi4iu6 & R0nhu6));
assign Xi4iu6 = (Shhpw6[6] & Iqzhu6);
assign Zevow6 = (~(Sevow6 & Kj6ju6));
assign HWDATA[5] = (~(Nfvow6 & Ufvow6));
assign Ufvow6 = (~(Oh4iu6 & R0nhu6));
assign Oh4iu6 = (Shhpw6[5] & Iqzhu6);
assign Nfvow6 = (~(Sevow6 & Eg6ju6));
assign HWDATA[4] = (~(Bgvow6 & Igvow6));
assign Igvow6 = (~(H34iu6 & R0nhu6));
assign H34iu6 = (Shhpw6[4] & Iqzhu6);
assign Bgvow6 = (~(Sevow6 & Zw4ju6));
assign HWDATA[3] = (~(Pgvow6 & Wgvow6));
assign Wgvow6 = (~(Df4iu6 & R0nhu6));
assign Df4iu6 = (Shhpw6[3] & Iqzhu6);
assign Pgvow6 = (~(Sevow6 & G36ju6));
assign HWDATA[31] = (~(Dhvow6 & Khvow6));
assign Khvow6 = (Rhvow6 & Yhvow6);
assign Yhvow6 = (~(Gdqow6 & Aioiu6));
assign Aioiu6 = (~(Fivow6 & Mivow6));
assign Mivow6 = (Tivow6 & Ajvow6);
assign Ajvow6 = (Hjvow6 & Ojvow6);
assign Ojvow6 = (~(vis_r11_o[31] & Ljqow6));
assign Hjvow6 = (Vjvow6 & Ckvow6);
assign Ckvow6 = (~(vis_r9_o[31] & Qiqow6));
assign Vjvow6 = (~(Fkfpw6[31] & Dfqow6));
assign Tivow6 = (Jkvow6 & Qkvow6);
assign Qkvow6 = (~(vis_r10_o[31] & Sjqow6));
assign Jkvow6 = (~(vis_psp_o[29] & Yfqow6));
assign Fivow6 = (Xkvow6 & Elvow6);
assign Elvow6 = (Llvow6 & Slvow6);
assign Slvow6 = (~(vis_r12_o[31] & Hhqow6));
assign Llvow6 = (Zlvow6 & Gmvow6);
assign Gmvow6 = (~(vis_msp_o[29] & Fgqow6));
assign Zlvow6 = (~(vis_r14_o[31] & Ahqow6));
assign Xkvow6 = (Bxzhu6 & Nmvow6);
assign Nmvow6 = (~(vis_r8_o[31] & Gkqow6));
assign Bxzhu6 = (Umvow6 & Bnvow6);
assign Bnvow6 = (Invow6 & Pnvow6);
assign Pnvow6 = (Wnvow6 & Dovow6);
assign Dovow6 = (~(vis_r2_o[31] & Dmqow6));
assign Wnvow6 = (~(vis_r6_o[31] & Kmqow6));
assign Invow6 = (Kovow6 & Rovow6);
assign Rovow6 = (~(vis_r5_o[31] & Fnqow6));
assign Kovow6 = (~(vis_r4_o[31] & Mnqow6));
assign Umvow6 = (Yovow6 & Fpvow6);
assign Fpvow6 = (Mpvow6 & Tpvow6);
assign Tpvow6 = (~(vis_r1_o[31] & Voqow6));
assign Mpvow6 = (~(vis_r0_o[31] & Cpqow6));
assign Yovow6 = (Aqvow6 & Hqvow6);
assign Hqvow6 = (~(vis_r3_o[31] & Xpqow6));
assign Aqvow6 = (~(vis_r7_o[31] & Eqqow6));
assign Rhvow6 = (~(R0nhu6 & Lm1iu6));
assign Lm1iu6 = (Shhpw6[31] & Iqzhu6);
assign Dhvow6 = (Oqvow6 & Vqvow6);
assign Vqvow6 = (~(K0row6 & W89ju6));
assign HWDATA[30] = (~(Crvow6 & Jrvow6));
assign Jrvow6 = (Qrvow6 & Xrvow6);
assign Xrvow6 = (~(Gdqow6 & T6liu6));
assign T6liu6 = (~(Esvow6 & Lsvow6));
assign Lsvow6 = (Ssvow6 & Zsvow6);
assign Zsvow6 = (Gtvow6 & Ntvow6);
assign Ntvow6 = (~(vis_r11_o[30] & Ljqow6));
assign Gtvow6 = (Utvow6 & Buvow6);
assign Buvow6 = (~(vis_r10_o[30] & Sjqow6));
assign Utvow6 = (~(vis_r9_o[30] & Qiqow6));
assign Ssvow6 = (Iuvow6 & Puvow6);
assign Puvow6 = (~(Fkfpw6[30] & Dfqow6));
assign Iuvow6 = (~(vis_r12_o[30] & Hhqow6));
assign Esvow6 = (Wuvow6 & Dvvow6);
assign Dvvow6 = (Kvvow6 & Rvvow6);
assign Rvvow6 = (~(vis_r14_o[30] & Ahqow6));
assign Kvvow6 = (Yvvow6 & Fwvow6);
assign Fwvow6 = (~(vis_psp_o[28] & Yfqow6));
assign Yvvow6 = (~(vis_r8_o[30] & Gkqow6));
assign Wuvow6 = (Ixzhu6 & Mwvow6);
assign Mwvow6 = (~(vis_msp_o[28] & Fgqow6));
assign Ixzhu6 = (Twvow6 & Axvow6);
assign Axvow6 = (Hxvow6 & Oxvow6);
assign Oxvow6 = (Vxvow6 & Cyvow6);
assign Cyvow6 = (~(vis_r0_o[30] & Cpqow6));
assign Vxvow6 = (~(vis_r2_o[30] & Dmqow6));
assign Hxvow6 = (Jyvow6 & Qyvow6);
assign Qyvow6 = (~(vis_r5_o[30] & Fnqow6));
assign Jyvow6 = (~(vis_r4_o[30] & Mnqow6));
assign Twvow6 = (Xyvow6 & Ezvow6);
assign Ezvow6 = (Lzvow6 & Szvow6);
assign Szvow6 = (~(vis_r7_o[30] & Eqqow6));
assign Lzvow6 = (~(vis_r3_o[30] & Xpqow6));
assign Xyvow6 = (Zzvow6 & G0wow6);
assign G0wow6 = (~(vis_r1_o[30] & Voqow6));
assign Zzvow6 = (~(vis_r6_o[30] & Kmqow6));
assign Qrvow6 = (Naliu6 | Qaxiu6);
assign Naliu6 = (!T94iu6);
assign T94iu6 = (Shhpw6[30] & Iqzhu6);
assign Crvow6 = (N0wow6 & U0wow6);
assign U0wow6 = (~(K0row6 & T39ju6));
assign HWDATA[2] = (~(B1wow6 & I1wow6));
assign I1wow6 = (~(Ud4iu6 & R0nhu6));
assign Ud4iu6 = (Shhpw6[2] & Iqzhu6);
assign B1wow6 = (~(Sevow6 & Ot5ju6));
assign HWDATA[28] = (~(P1wow6 & W1wow6));
assign W1wow6 = (D2wow6 & K2wow6);
assign K2wow6 = (~(Gdqow6 & Po7ju6));
assign Po7ju6 = (~(R2wow6 & Y2wow6));
assign Y2wow6 = (F3wow6 & M3wow6);
assign M3wow6 = (T3wow6 & A4wow6);
assign A4wow6 = (~(vis_r11_o[28] & Ljqow6));
assign T3wow6 = (H4wow6 & O4wow6);
assign O4wow6 = (~(vis_r10_o[28] & Sjqow6));
assign H4wow6 = (~(vis_r9_o[28] & Qiqow6));
assign F3wow6 = (V4wow6 & C5wow6);
assign C5wow6 = (~(Fkfpw6[28] & Dfqow6));
assign V4wow6 = (~(vis_r12_o[28] & Hhqow6));
assign R2wow6 = (J5wow6 & Q5wow6);
assign Q5wow6 = (X5wow6 & E6wow6);
assign E6wow6 = (~(vis_r14_o[28] & Ahqow6));
assign X5wow6 = (L6wow6 & S6wow6);
assign S6wow6 = (~(vis_psp_o[26] & Yfqow6));
assign L6wow6 = (~(vis_r8_o[28] & Gkqow6));
assign J5wow6 = (Dyzhu6 & Z6wow6);
assign Z6wow6 = (~(vis_msp_o[26] & Fgqow6));
assign Dyzhu6 = (G7wow6 & N7wow6);
assign N7wow6 = (U7wow6 & B8wow6);
assign B8wow6 = (I8wow6 & P8wow6);
assign P8wow6 = (~(vis_r0_o[28] & Cpqow6));
assign I8wow6 = (~(vis_r2_o[28] & Dmqow6));
assign U7wow6 = (W8wow6 & D9wow6);
assign D9wow6 = (~(vis_r5_o[28] & Fnqow6));
assign W8wow6 = (~(vis_r4_o[28] & Mnqow6));
assign G7wow6 = (K9wow6 & R9wow6);
assign R9wow6 = (Y9wow6 & Fawow6);
assign Fawow6 = (~(vis_r7_o[28] & Eqqow6));
assign Y9wow6 = (~(vis_r3_o[28] & Xpqow6));
assign K9wow6 = (Mawow6 & Tawow6);
assign Tawow6 = (~(vis_r1_o[28] & Voqow6));
assign Mawow6 = (~(vis_r6_o[28] & Kmqow6));
assign D2wow6 = (Zeniu6 | Qaxiu6);
assign Zeniu6 = (!F94iu6);
assign F94iu6 = (Shhpw6[28] & Iqzhu6);
assign P1wow6 = (Abwow6 & Hbwow6);
assign Hbwow6 = (~(K0row6 & Rv8ju6));
assign HWDATA[27] = (~(Obwow6 & Vbwow6));
assign Vbwow6 = (Ccwow6 & Jcwow6);
assign Jcwow6 = (~(Gdqow6 & A67ju6));
assign A67ju6 = (~(Qcwow6 & Xcwow6));
assign Xcwow6 = (Edwow6 & Ldwow6);
assign Ldwow6 = (Sdwow6 & Zdwow6);
assign Zdwow6 = (~(Fkfpw6[27] & Dfqow6));
assign Sdwow6 = (Gewow6 & Newow6);
assign Newow6 = (~(vis_psp_o[25] & Yfqow6));
assign Gewow6 = (~(vis_msp_o[25] & Fgqow6));
assign Edwow6 = (Uewow6 & Bfwow6);
assign Bfwow6 = (~(vis_r14_o[27] & Ahqow6));
assign Uewow6 = (~(vis_r12_o[27] & Hhqow6));
assign Qcwow6 = (Ifwow6 & Pfwow6);
assign Pfwow6 = (Wfwow6 & Dgwow6);
assign Dgwow6 = (~(vis_r9_o[27] & Qiqow6));
assign Wfwow6 = (Kgwow6 & Rgwow6);
assign Rgwow6 = (~(vis_r11_o[27] & Ljqow6));
assign Kgwow6 = (~(vis_r10_o[27] & Sjqow6));
assign Ifwow6 = (Kyzhu6 & Ygwow6);
assign Ygwow6 = (~(vis_r8_o[27] & Gkqow6));
assign Kyzhu6 = (Fhwow6 & Mhwow6);
assign Mhwow6 = (Thwow6 & Aiwow6);
assign Aiwow6 = (Hiwow6 & Oiwow6);
assign Oiwow6 = (~(vis_r2_o[27] & Dmqow6));
assign Hiwow6 = (~(vis_r6_o[27] & Kmqow6));
assign Thwow6 = (Viwow6 & Cjwow6);
assign Cjwow6 = (~(vis_r5_o[27] & Fnqow6));
assign Viwow6 = (~(vis_r4_o[27] & Mnqow6));
assign Fhwow6 = (Jjwow6 & Qjwow6);
assign Qjwow6 = (Xjwow6 & Ekwow6);
assign Ekwow6 = (~(vis_r1_o[27] & Voqow6));
assign Xjwow6 = (~(vis_r0_o[27] & Cpqow6));
assign Jjwow6 = (Lkwow6 & Skwow6);
assign Skwow6 = (~(vis_r3_o[27] & Xpqow6));
assign Lkwow6 = (~(vis_r7_o[27] & Eqqow6));
assign Ccwow6 = (U3liu6 | Qaxiu6);
assign U3liu6 = (!Y84iu6);
assign Y84iu6 = (Shhpw6[27] & Iqzhu6);
assign Obwow6 = (Zkwow6 & Glwow6);
assign Glwow6 = (~(K0row6 & In8ju6));
assign K0row6 = (!Nlwow6);
assign HWDATA[26] = (~(Ulwow6 & Bmwow6));
assign Bmwow6 = (Imwow6 & Pmwow6);
assign Pmwow6 = (~(Gdqow6 & Z17ju6));
assign Z17ju6 = (~(Wmwow6 & Dnwow6));
assign Dnwow6 = (Knwow6 & Rnwow6);
assign Rnwow6 = (Ynwow6 & Fowow6);
assign Fowow6 = (~(Fkfpw6[26] & Dfqow6));
assign Ynwow6 = (Mowow6 & Towow6);
assign Towow6 = (~(vis_psp_o[24] & Yfqow6));
assign Mowow6 = (~(vis_msp_o[24] & Fgqow6));
assign Knwow6 = (Apwow6 & Hpwow6);
assign Hpwow6 = (~(vis_r14_o[26] & Ahqow6));
assign Apwow6 = (~(vis_r12_o[26] & Hhqow6));
assign Wmwow6 = (Opwow6 & Vpwow6);
assign Vpwow6 = (Cqwow6 & Jqwow6);
assign Jqwow6 = (~(vis_r9_o[26] & Qiqow6));
assign Cqwow6 = (Qqwow6 & Xqwow6);
assign Xqwow6 = (~(vis_r11_o[26] & Ljqow6));
assign Qqwow6 = (~(vis_r10_o[26] & Sjqow6));
assign Opwow6 = (Ryzhu6 & Erwow6);
assign Erwow6 = (~(vis_r8_o[26] & Gkqow6));
assign Ryzhu6 = (Lrwow6 & Srwow6);
assign Srwow6 = (Zrwow6 & Gswow6);
assign Gswow6 = (Nswow6 & Uswow6);
assign Uswow6 = (~(vis_r2_o[26] & Dmqow6));
assign Nswow6 = (~(vis_r6_o[26] & Kmqow6));
assign Zrwow6 = (Btwow6 & Itwow6);
assign Itwow6 = (~(vis_r5_o[26] & Fnqow6));
assign Btwow6 = (~(vis_r4_o[26] & Mnqow6));
assign Lrwow6 = (Ptwow6 & Wtwow6);
assign Wtwow6 = (Duwow6 & Kuwow6);
assign Kuwow6 = (~(vis_r1_o[26] & Voqow6));
assign Duwow6 = (~(vis_r0_o[26] & Cpqow6));
assign Ptwow6 = (Ruwow6 & Yuwow6);
assign Yuwow6 = (~(vis_r3_o[26] & Xpqow6));
assign Ruwow6 = (~(vis_r7_o[26] & Eqqow6));
assign Imwow6 = (C1liu6 | Qaxiu6);
assign C1liu6 = (!R84iu6);
assign R84iu6 = (Shhpw6[26] & Iqzhu6);
assign Ulwow6 = (Fvwow6 & Mvwow6);
assign Mvwow6 = (Nlwow6 | Ka8ju6);
assign HWDATA[25] = (~(Tvwow6 & Awwow6));
assign Awwow6 = (Hwwow6 & Owwow6);
assign Owwow6 = (Nlwow6 | I28ju6);
assign I28ju6 = (Vwwow6 & Cxwow6);
assign Cxwow6 = (Jxwow6 & Qxwow6);
assign Qxwow6 = (Xxwow6 & Eywow6);
assign Eywow6 = (~(vis_r11_o[9] & Ljqow6));
assign Xxwow6 = (Lywow6 & Sywow6);
assign Sywow6 = (~(vis_r10_o[9] & Sjqow6));
assign Lywow6 = (~(vis_r9_o[9] & Qiqow6));
assign Jxwow6 = (Zywow6 & Gzwow6);
assign Gzwow6 = (~(Fkfpw6[9] & Dfqow6));
assign Zywow6 = (~(vis_r12_o[9] & Hhqow6));
assign Vwwow6 = (Nzwow6 & Uzwow6);
assign Uzwow6 = (B0xow6 & I0xow6);
assign I0xow6 = (~(vis_r14_o[9] & Ahqow6));
assign B0xow6 = (P0xow6 & W0xow6);
assign W0xow6 = (~(vis_psp_o[7] & Yfqow6));
assign P0xow6 = (~(vis_r8_o[9] & Gkqow6));
assign Nzwow6 = (Evzhu6 & D1xow6);
assign D1xow6 = (~(vis_msp_o[7] & Fgqow6));
assign Evzhu6 = (K1xow6 & R1xow6);
assign R1xow6 = (Y1xow6 & F2xow6);
assign F2xow6 = (M2xow6 & T2xow6);
assign T2xow6 = (~(vis_r0_o[9] & Cpqow6));
assign M2xow6 = (~(vis_r2_o[9] & Dmqow6));
assign Y1xow6 = (A3xow6 & H3xow6);
assign H3xow6 = (~(vis_r5_o[9] & Fnqow6));
assign A3xow6 = (~(vis_r4_o[9] & Mnqow6));
assign K1xow6 = (O3xow6 & V3xow6);
assign V3xow6 = (C4xow6 & J4xow6);
assign J4xow6 = (~(vis_r7_o[9] & Eqqow6));
assign C4xow6 = (~(vis_r3_o[9] & Xpqow6));
assign O3xow6 = (Q4xow6 & X4xow6);
assign X4xow6 = (~(vis_r1_o[9] & Voqow6));
assign Q4xow6 = (~(vis_r6_o[9] & Kmqow6));
assign Hwwow6 = (~(Gdqow6 & Goliu6));
assign Goliu6 = (~(E5xow6 & L5xow6));
assign L5xow6 = (S5xow6 & Z5xow6);
assign Z5xow6 = (G6xow6 & N6xow6);
assign N6xow6 = (~(Fkfpw6[25] & Dfqow6));
assign G6xow6 = (U6xow6 & B7xow6);
assign B7xow6 = (~(vis_psp_o[23] & Yfqow6));
assign U6xow6 = (~(vis_msp_o[23] & Fgqow6));
assign S5xow6 = (I7xow6 & P7xow6);
assign P7xow6 = (~(vis_r14_o[25] & Ahqow6));
assign I7xow6 = (~(vis_r12_o[25] & Hhqow6));
assign E5xow6 = (W7xow6 & D8xow6);
assign D8xow6 = (K8xow6 & R8xow6);
assign R8xow6 = (~(vis_r9_o[25] & Qiqow6));
assign K8xow6 = (Y8xow6 & F9xow6);
assign F9xow6 = (~(vis_r11_o[25] & Ljqow6));
assign Y8xow6 = (~(vis_r10_o[25] & Sjqow6));
assign W7xow6 = (Yyzhu6 & M9xow6);
assign M9xow6 = (~(vis_r8_o[25] & Gkqow6));
assign Yyzhu6 = (T9xow6 & Aaxow6);
assign Aaxow6 = (Haxow6 & Oaxow6);
assign Oaxow6 = (Vaxow6 & Cbxow6);
assign Cbxow6 = (~(vis_r2_o[25] & Dmqow6));
assign Vaxow6 = (~(vis_r6_o[25] & Kmqow6));
assign Haxow6 = (Jbxow6 & Qbxow6);
assign Qbxow6 = (~(vis_r5_o[25] & Fnqow6));
assign Jbxow6 = (~(vis_r4_o[25] & Mnqow6));
assign T9xow6 = (Xbxow6 & Ecxow6);
assign Ecxow6 = (Lcxow6 & Scxow6);
assign Scxow6 = (~(vis_r1_o[25] & Voqow6));
assign Lcxow6 = (~(vis_r0_o[25] & Cpqow6));
assign Xbxow6 = (Zcxow6 & Gdxow6);
assign Gdxow6 = (~(vis_r3_o[25] & Xpqow6));
assign Zcxow6 = (~(vis_r7_o[25] & Eqqow6));
assign Tvwow6 = (Acvow6 & Ndxow6);
assign Ndxow6 = (Asliu6 | Qaxiu6);
assign Asliu6 = (!K84iu6);
assign K84iu6 = (Shhpw6[25] & Iqzhu6);
assign Acvow6 = (~(Udxow6 & Znliu6));
assign HWDATA[24] = (~(Bexow6 & Iexow6));
assign Iexow6 = (Pexow6 & Wexow6);
assign Wexow6 = (Nlwow6 | Cz7ju6);
assign Cz7ju6 = (Dfxow6 & Kfxow6);
assign Kfxow6 = (Rfxow6 & Yfxow6);
assign Yfxow6 = (Fgxow6 & Mgxow6);
assign Mgxow6 = (~(vis_r11_o[8] & Ljqow6));
assign Fgxow6 = (Tgxow6 & Ahxow6);
assign Ahxow6 = (~(vis_r9_o[8] & Qiqow6));
assign Tgxow6 = (~(Fkfpw6[8] & Dfqow6));
assign Rfxow6 = (Hhxow6 & Ohxow6);
assign Ohxow6 = (~(vis_r10_o[8] & Sjqow6));
assign Hhxow6 = (~(vis_psp_o[6] & Yfqow6));
assign Dfxow6 = (Vhxow6 & Cixow6);
assign Cixow6 = (Jixow6 & Qixow6);
assign Qixow6 = (~(vis_r12_o[8] & Hhqow6));
assign Jixow6 = (Xixow6 & Ejxow6);
assign Ejxow6 = (~(vis_msp_o[6] & Fgqow6));
assign Xixow6 = (~(vis_r14_o[8] & Ahqow6));
assign Vhxow6 = (Lvzhu6 & Ljxow6);
assign Ljxow6 = (~(vis_r8_o[8] & Gkqow6));
assign Lvzhu6 = (Sjxow6 & Zjxow6);
assign Zjxow6 = (Gkxow6 & Nkxow6);
assign Nkxow6 = (Ukxow6 & Blxow6);
assign Blxow6 = (~(vis_r2_o[8] & Dmqow6));
assign Ukxow6 = (~(vis_r6_o[8] & Kmqow6));
assign Gkxow6 = (Ilxow6 & Plxow6);
assign Plxow6 = (~(vis_r5_o[8] & Fnqow6));
assign Ilxow6 = (~(vis_r4_o[8] & Mnqow6));
assign Sjxow6 = (Wlxow6 & Dmxow6);
assign Dmxow6 = (Kmxow6 & Rmxow6);
assign Rmxow6 = (~(vis_r1_o[8] & Voqow6));
assign Kmxow6 = (~(vis_r0_o[8] & Cpqow6));
assign Wlxow6 = (Ymxow6 & Fnxow6);
assign Fnxow6 = (~(vis_r3_o[8] & Xpqow6));
assign Ymxow6 = (~(vis_r7_o[8] & Eqqow6));
assign Nlwow6 = (~(Mnxow6 & Sevow6));
assign Pexow6 = (~(Gdqow6 & Fy6ju6));
assign Fy6ju6 = (~(Tnxow6 & Aoxow6));
assign Aoxow6 = (Hoxow6 & Ooxow6);
assign Ooxow6 = (Voxow6 & Cpxow6);
assign Cpxow6 = (~(Fkfpw6[24] & Dfqow6));
assign Voxow6 = (Jpxow6 & Qpxow6);
assign Qpxow6 = (~(vis_psp_o[22] & Yfqow6));
assign Jpxow6 = (~(vis_msp_o[22] & Fgqow6));
assign Hoxow6 = (Xpxow6 & Eqxow6);
assign Eqxow6 = (~(vis_r14_o[24] & Ahqow6));
assign Xpxow6 = (~(vis_r12_o[24] & Hhqow6));
assign Tnxow6 = (Lqxow6 & Sqxow6);
assign Sqxow6 = (Zqxow6 & Grxow6);
assign Grxow6 = (~(vis_r9_o[24] & Qiqow6));
assign Zqxow6 = (Nrxow6 & Urxow6);
assign Urxow6 = (~(vis_r11_o[24] & Ljqow6));
assign Nrxow6 = (~(vis_r10_o[24] & Sjqow6));
assign Lqxow6 = (Fzzhu6 & Bsxow6);
assign Bsxow6 = (~(vis_r8_o[24] & Gkqow6));
assign Fzzhu6 = (Isxow6 & Psxow6);
assign Psxow6 = (Wsxow6 & Dtxow6);
assign Dtxow6 = (Ktxow6 & Rtxow6);
assign Rtxow6 = (~(vis_r2_o[24] & Dmqow6));
assign Ktxow6 = (~(vis_r6_o[24] & Kmqow6));
assign Wsxow6 = (Ytxow6 & Fuxow6);
assign Fuxow6 = (~(vis_r5_o[24] & Fnqow6));
assign Ytxow6 = (~(vis_r4_o[24] & Mnqow6));
assign Isxow6 = (Muxow6 & Tuxow6);
assign Tuxow6 = (Avxow6 & Hvxow6);
assign Hvxow6 = (~(vis_r1_o[24] & Voqow6));
assign Avxow6 = (~(vis_r0_o[24] & Cpqow6));
assign Muxow6 = (Ovxow6 & Vvxow6);
assign Vvxow6 = (~(vis_r3_o[24] & Xpqow6));
assign Ovxow6 = (~(vis_r7_o[24] & Eqqow6));
assign Bexow6 = (Jdvow6 & Cwxow6);
assign Cwxow6 = (Rykiu6 | Qaxiu6);
assign Rykiu6 = (!D84iu6);
assign D84iu6 = (Shhpw6[24] & Iqzhu6);
assign Jdvow6 = (~(Udxow6 & L35ju6));
assign HWDATA[23] = (~(Jwxow6 & Qwxow6));
assign Qwxow6 = (~(Lcqow6 & Uo6ju6));
assign Jwxow6 = (Xwxow6 & Exxow6);
assign Exxow6 = (Ox9iu6 | Qaxiu6);
assign Ox9iu6 = (!W74iu6);
assign W74iu6 = (Shhpw6[23] & Iqzhu6);
assign Xwxow6 = (~(Gdqow6 & Xg5ju6));
assign Xg5ju6 = (~(Lxxow6 & Sxxow6));
assign Sxxow6 = (Zxxow6 & Gyxow6);
assign Gyxow6 = (Nyxow6 & Uyxow6);
assign Uyxow6 = (~(Fkfpw6[23] & Dfqow6));
assign Nyxow6 = (Bzxow6 & Izxow6);
assign Izxow6 = (~(vis_psp_o[21] & Yfqow6));
assign Bzxow6 = (~(vis_msp_o[21] & Fgqow6));
assign Zxxow6 = (Pzxow6 & Wzxow6);
assign Wzxow6 = (~(vis_r14_o[23] & Ahqow6));
assign Pzxow6 = (~(vis_r12_o[23] & Hhqow6));
assign Lxxow6 = (D0yow6 & K0yow6);
assign K0yow6 = (R0yow6 & Y0yow6);
assign Y0yow6 = (~(vis_r9_o[23] & Qiqow6));
assign R0yow6 = (F1yow6 & M1yow6);
assign M1yow6 = (~(vis_r11_o[23] & Ljqow6));
assign F1yow6 = (~(vis_r10_o[23] & Sjqow6));
assign D0yow6 = (Mzzhu6 & T1yow6);
assign T1yow6 = (~(vis_r8_o[23] & Gkqow6));
assign Mzzhu6 = (A2yow6 & H2yow6);
assign H2yow6 = (O2yow6 & V2yow6);
assign V2yow6 = (C3yow6 & J3yow6);
assign J3yow6 = (~(vis_r2_o[23] & Dmqow6));
assign C3yow6 = (~(vis_r6_o[23] & Kmqow6));
assign O2yow6 = (Q3yow6 & X3yow6);
assign X3yow6 = (~(vis_r5_o[23] & Fnqow6));
assign Q3yow6 = (~(vis_r4_o[23] & Mnqow6));
assign A2yow6 = (E4yow6 & L4yow6);
assign L4yow6 = (S4yow6 & Z4yow6);
assign Z4yow6 = (~(vis_r1_o[23] & Voqow6));
assign S4yow6 = (~(vis_r0_o[23] & Cpqow6));
assign E4yow6 = (G5yow6 & N5yow6);
assign N5yow6 = (~(vis_r3_o[23] & Xpqow6));
assign G5yow6 = (~(vis_r7_o[23] & Eqqow6));
assign HWDATA[22] = (~(U5yow6 & B6yow6));
assign B6yow6 = (~(Lcqow6 & Kj6ju6));
assign U5yow6 = (I6yow6 & P6yow6);
assign P6yow6 = (~(P74iu6 & R0nhu6));
assign P74iu6 = (Shhpw6[22] & Iqzhu6);
assign I6yow6 = (~(Gdqow6 & V3aju6));
assign V3aju6 = (~(W6yow6 & D7yow6));
assign D7yow6 = (K7yow6 & R7yow6);
assign R7yow6 = (Y7yow6 & F8yow6);
assign F8yow6 = (~(Fkfpw6[22] & Dfqow6));
assign Y7yow6 = (M8yow6 & T8yow6);
assign T8yow6 = (~(vis_psp_o[20] & Yfqow6));
assign M8yow6 = (~(vis_msp_o[20] & Fgqow6));
assign K7yow6 = (A9yow6 & H9yow6);
assign H9yow6 = (~(vis_r14_o[22] & Ahqow6));
assign A9yow6 = (~(vis_r12_o[22] & Hhqow6));
assign W6yow6 = (O9yow6 & V9yow6);
assign V9yow6 = (Cayow6 & Jayow6);
assign Jayow6 = (~(vis_r9_o[22] & Qiqow6));
assign Cayow6 = (Qayow6 & Xayow6);
assign Xayow6 = (~(vis_r11_o[22] & Ljqow6));
assign Qayow6 = (~(vis_r10_o[22] & Sjqow6));
assign O9yow6 = (Tzzhu6 & Ebyow6);
assign Ebyow6 = (~(vis_r8_o[22] & Gkqow6));
assign Tzzhu6 = (Lbyow6 & Sbyow6);
assign Sbyow6 = (Zbyow6 & Gcyow6);
assign Gcyow6 = (Ncyow6 & Ucyow6);
assign Ucyow6 = (~(vis_r2_o[22] & Dmqow6));
assign Ncyow6 = (~(vis_r6_o[22] & Kmqow6));
assign Zbyow6 = (Bdyow6 & Idyow6);
assign Idyow6 = (~(vis_r5_o[22] & Fnqow6));
assign Bdyow6 = (~(vis_r4_o[22] & Mnqow6));
assign Lbyow6 = (Pdyow6 & Wdyow6);
assign Wdyow6 = (Deyow6 & Keyow6);
assign Keyow6 = (~(vis_r1_o[22] & Voqow6));
assign Deyow6 = (~(vis_r0_o[22] & Cpqow6));
assign Pdyow6 = (Reyow6 & Yeyow6);
assign Yeyow6 = (~(vis_r3_o[22] & Xpqow6));
assign Reyow6 = (~(vis_r7_o[22] & Eqqow6));
assign HWDATA[21] = (~(Ffyow6 & Mfyow6));
assign Mfyow6 = (~(Lcqow6 & Eg6ju6));
assign Ffyow6 = (Tfyow6 & Agyow6);
assign Agyow6 = (Yxliu6 | Qaxiu6);
assign Yxliu6 = (!I74iu6);
assign I74iu6 = (Shhpw6[21] & Iqzhu6);
assign Tfyow6 = (~(Gdqow6 & Xx9ju6));
assign Xx9ju6 = (~(Hgyow6 & Ogyow6));
assign Ogyow6 = (Vgyow6 & Chyow6);
assign Chyow6 = (Jhyow6 & Qhyow6);
assign Qhyow6 = (~(Fkfpw6[21] & Dfqow6));
assign Jhyow6 = (Xhyow6 & Eiyow6);
assign Eiyow6 = (~(vis_psp_o[19] & Yfqow6));
assign Xhyow6 = (~(vis_msp_o[19] & Fgqow6));
assign Vgyow6 = (Liyow6 & Siyow6);
assign Siyow6 = (~(vis_r14_o[21] & Ahqow6));
assign Liyow6 = (~(vis_r12_o[21] & Hhqow6));
assign Hgyow6 = (Ziyow6 & Gjyow6);
assign Gjyow6 = (Njyow6 & Ujyow6);
assign Ujyow6 = (~(vis_r9_o[21] & Qiqow6));
assign Njyow6 = (Bkyow6 & Ikyow6);
assign Ikyow6 = (~(vis_r11_o[21] & Ljqow6));
assign Bkyow6 = (~(vis_r10_o[21] & Sjqow6));
assign Ziyow6 = (A00iu6 & Pkyow6);
assign Pkyow6 = (~(vis_r8_o[21] & Gkqow6));
assign A00iu6 = (Wkyow6 & Dlyow6);
assign Dlyow6 = (Klyow6 & Rlyow6);
assign Rlyow6 = (Ylyow6 & Fmyow6);
assign Fmyow6 = (~(vis_r2_o[21] & Dmqow6));
assign Ylyow6 = (~(vis_r6_o[21] & Kmqow6));
assign Klyow6 = (Mmyow6 & Tmyow6);
assign Tmyow6 = (~(vis_r5_o[21] & Fnqow6));
assign Mmyow6 = (~(vis_r4_o[21] & Mnqow6));
assign Wkyow6 = (Anyow6 & Hnyow6);
assign Hnyow6 = (Onyow6 & Vnyow6);
assign Vnyow6 = (~(vis_r1_o[21] & Voqow6));
assign Onyow6 = (~(vis_r0_o[21] & Cpqow6));
assign Anyow6 = (Coyow6 & Joyow6);
assign Joyow6 = (~(vis_r3_o[21] & Xpqow6));
assign Coyow6 = (~(vis_r7_o[21] & Eqqow6));
assign HWDATA[20] = (~(Qoyow6 & Xoyow6));
assign Xoyow6 = (~(Lcqow6 & Zw4ju6));
assign Qoyow6 = (Epyow6 & Lpyow6);
assign Lpyow6 = (~(B74iu6 & R0nhu6));
assign B74iu6 = (Shhpw6[20] & Iqzhu6);
assign Epyow6 = (~(Gdqow6 & Wt9ju6));
assign Wt9ju6 = (~(Spyow6 & Zpyow6));
assign Zpyow6 = (Gqyow6 & Nqyow6);
assign Nqyow6 = (Uqyow6 & Bryow6);
assign Bryow6 = (~(Fkfpw6[20] & Dfqow6));
assign Uqyow6 = (Iryow6 & Pryow6);
assign Pryow6 = (~(vis_psp_o[18] & Yfqow6));
assign Iryow6 = (~(vis_msp_o[18] & Fgqow6));
assign Gqyow6 = (Wryow6 & Dsyow6);
assign Dsyow6 = (~(vis_r14_o[20] & Ahqow6));
assign Wryow6 = (~(vis_r12_o[20] & Hhqow6));
assign Spyow6 = (Ksyow6 & Rsyow6);
assign Rsyow6 = (Ysyow6 & Ftyow6);
assign Ftyow6 = (~(vis_r9_o[20] & Qiqow6));
assign Ysyow6 = (Mtyow6 & Ttyow6);
assign Ttyow6 = (~(vis_r11_o[20] & Ljqow6));
assign Mtyow6 = (~(vis_r10_o[20] & Sjqow6));
assign Ksyow6 = (H00iu6 & Auyow6);
assign Auyow6 = (~(vis_r8_o[20] & Gkqow6));
assign H00iu6 = (Huyow6 & Ouyow6);
assign Ouyow6 = (Vuyow6 & Cvyow6);
assign Cvyow6 = (Jvyow6 & Qvyow6);
assign Qvyow6 = (~(vis_r2_o[20] & Dmqow6));
assign Jvyow6 = (~(vis_r6_o[20] & Kmqow6));
assign Vuyow6 = (Xvyow6 & Ewyow6);
assign Ewyow6 = (~(vis_r5_o[20] & Fnqow6));
assign Xvyow6 = (~(vis_r4_o[20] & Mnqow6));
assign Huyow6 = (Lwyow6 & Swyow6);
assign Swyow6 = (Zwyow6 & Gxyow6);
assign Gxyow6 = (~(vis_r1_o[20] & Voqow6));
assign Zwyow6 = (~(vis_r0_o[20] & Cpqow6));
assign Lwyow6 = (Nxyow6 & Uxyow6);
assign Uxyow6 = (~(vis_r3_o[20] & Xpqow6));
assign Nxyow6 = (~(vis_r7_o[20] & Eqqow6));
assign HWDATA[1] = (~(Byyow6 & Iyyow6));
assign Iyyow6 = (A34iu6 | Qaxiu6);
assign A34iu6 = (!O34iu6);
assign O34iu6 = (Shhpw6[1] & Iqzhu6);
assign Byyow6 = (~(Sevow6 & Znliu6));
assign HWDATA[19] = (~(Pyyow6 & Wyyow6));
assign Wyyow6 = (~(Lcqow6 & G36ju6));
assign Pyyow6 = (Dzyow6 & Kzyow6);
assign Kzyow6 = (~(U64iu6 & R0nhu6));
assign U64iu6 = (Shhpw6[19] & Iqzhu6);
assign Dzyow6 = (~(Gdqow6 & Vp9ju6));
assign Vp9ju6 = (~(Rzyow6 & Yzyow6));
assign Yzyow6 = (F0zow6 & M0zow6);
assign M0zow6 = (T0zow6 & A1zow6);
assign A1zow6 = (~(Fkfpw6[19] & Dfqow6));
assign T0zow6 = (H1zow6 & O1zow6);
assign O1zow6 = (~(vis_psp_o[17] & Yfqow6));
assign H1zow6 = (~(vis_msp_o[17] & Fgqow6));
assign F0zow6 = (V1zow6 & C2zow6);
assign C2zow6 = (~(vis_r14_o[19] & Ahqow6));
assign V1zow6 = (~(vis_r12_o[19] & Hhqow6));
assign Rzyow6 = (J2zow6 & Q2zow6);
assign Q2zow6 = (X2zow6 & E3zow6);
assign E3zow6 = (~(vis_r9_o[19] & Qiqow6));
assign X2zow6 = (L3zow6 & S3zow6);
assign S3zow6 = (~(vis_r11_o[19] & Ljqow6));
assign L3zow6 = (~(vis_r10_o[19] & Sjqow6));
assign J2zow6 = (V00iu6 & Z3zow6);
assign Z3zow6 = (~(vis_r8_o[19] & Gkqow6));
assign V00iu6 = (G4zow6 & N4zow6);
assign N4zow6 = (U4zow6 & B5zow6);
assign B5zow6 = (I5zow6 & P5zow6);
assign P5zow6 = (~(vis_r2_o[19] & Dmqow6));
assign I5zow6 = (~(vis_r6_o[19] & Kmqow6));
assign U4zow6 = (W5zow6 & D6zow6);
assign D6zow6 = (~(vis_r5_o[19] & Fnqow6));
assign W5zow6 = (~(vis_r4_o[19] & Mnqow6));
assign G4zow6 = (K6zow6 & R6zow6);
assign R6zow6 = (Y6zow6 & F7zow6);
assign F7zow6 = (~(vis_r1_o[19] & Voqow6));
assign Y6zow6 = (~(vis_r0_o[19] & Cpqow6));
assign K6zow6 = (M7zow6 & T7zow6);
assign T7zow6 = (~(vis_r3_o[19] & Xpqow6));
assign M7zow6 = (~(vis_r7_o[19] & Eqqow6));
assign HWDATA[18] = (~(A8zow6 & H8zow6));
assign H8zow6 = (~(Lcqow6 & Ot5ju6));
assign A8zow6 = (O8zow6 & V8zow6);
assign V8zow6 = (~(N64iu6 & R0nhu6));
assign N64iu6 = (Shhpw6[18] & Iqzhu6);
assign O8zow6 = (~(Gdqow6 & Gl9ju6));
assign Gl9ju6 = (~(C9zow6 & J9zow6));
assign J9zow6 = (Q9zow6 & X9zow6);
assign X9zow6 = (Eazow6 & Lazow6);
assign Lazow6 = (~(Fkfpw6[18] & Dfqow6));
assign Eazow6 = (Sazow6 & Zazow6);
assign Zazow6 = (~(vis_psp_o[16] & Yfqow6));
assign Sazow6 = (~(vis_msp_o[16] & Fgqow6));
assign Q9zow6 = (Gbzow6 & Nbzow6);
assign Nbzow6 = (~(vis_r14_o[18] & Ahqow6));
assign Gbzow6 = (~(vis_r12_o[18] & Hhqow6));
assign C9zow6 = (Ubzow6 & Bczow6);
assign Bczow6 = (Iczow6 & Pczow6);
assign Pczow6 = (~(vis_r9_o[18] & Qiqow6));
assign Iczow6 = (Wczow6 & Ddzow6);
assign Ddzow6 = (~(vis_r11_o[18] & Ljqow6));
assign Wczow6 = (~(vis_r10_o[18] & Sjqow6));
assign Ubzow6 = (C10iu6 & Kdzow6);
assign Kdzow6 = (~(vis_r8_o[18] & Gkqow6));
assign C10iu6 = (Rdzow6 & Ydzow6);
assign Ydzow6 = (Fezow6 & Mezow6);
assign Mezow6 = (Tezow6 & Afzow6);
assign Afzow6 = (~(vis_r2_o[18] & Dmqow6));
assign Tezow6 = (~(vis_r6_o[18] & Kmqow6));
assign Fezow6 = (Hfzow6 & Ofzow6);
assign Ofzow6 = (~(vis_r5_o[18] & Fnqow6));
assign Hfzow6 = (~(vis_r4_o[18] & Mnqow6));
assign Rdzow6 = (Vfzow6 & Cgzow6);
assign Cgzow6 = (Jgzow6 & Qgzow6);
assign Qgzow6 = (~(vis_r1_o[18] & Voqow6));
assign Jgzow6 = (~(vis_r0_o[18] & Cpqow6));
assign Vfzow6 = (Xgzow6 & Ehzow6);
assign Ehzow6 = (~(vis_r3_o[18] & Xpqow6));
assign Xgzow6 = (~(vis_r7_o[18] & Eqqow6));
assign HWDATA[17] = (~(Lhzow6 & Shzow6));
assign Shzow6 = (~(Lcqow6 & Znliu6));
assign Znliu6 = (~(Zhzow6 & Gizow6));
assign Gizow6 = (Nizow6 & Uizow6);
assign Uizow6 = (Bjzow6 & Ijzow6);
assign Ijzow6 = (~(Fkfpw6[1] & Dfqow6));
assign Bjzow6 = (~(vis_r14_o[1] & Ahqow6));
assign Nizow6 = (Pjzow6 & Wjzow6);
assign Wjzow6 = (~(vis_r12_o[1] & Hhqow6));
assign Pjzow6 = (~(vis_r11_o[1] & Ljqow6));
assign Zhzow6 = (Dkzow6 & Kkzow6);
assign Kkzow6 = (Rkzow6 & Ykzow6);
assign Ykzow6 = (~(vis_r10_o[1] & Sjqow6));
assign Rkzow6 = (~(vis_r9_o[1] & Qiqow6));
assign Dkzow6 = (O00iu6 & Flzow6);
assign Flzow6 = (~(vis_r8_o[1] & Gkqow6));
assign O00iu6 = (Mlzow6 & Tlzow6);
assign Tlzow6 = (Amzow6 & Hmzow6);
assign Hmzow6 = (Omzow6 & Vmzow6);
assign Vmzow6 = (~(vis_r0_o[1] & Cpqow6));
assign Omzow6 = (~(vis_r2_o[1] & Dmqow6));
assign Amzow6 = (Cnzow6 & Jnzow6);
assign Jnzow6 = (~(vis_r5_o[1] & Fnqow6));
assign Cnzow6 = (~(vis_r4_o[1] & Mnqow6));
assign Mlzow6 = (Qnzow6 & Xnzow6);
assign Xnzow6 = (Eozow6 & Lozow6);
assign Lozow6 = (~(vis_r7_o[1] & Eqqow6));
assign Eozow6 = (~(vis_r3_o[1] & Xpqow6));
assign Qnzow6 = (Sozow6 & Zozow6);
assign Zozow6 = (~(vis_r1_o[1] & Voqow6));
assign Sozow6 = (~(vis_r6_o[1] & Kmqow6));
assign Lcqow6 = (Gpzow6 & Qaxiu6);
assign Gpzow6 = (~(L3ehu6 & X71iu6));
assign Lhzow6 = (Npzow6 & Upzow6);
assign Upzow6 = (~(Gdqow6 & Fh9ju6));
assign Fh9ju6 = (~(Bqzow6 & Iqzow6));
assign Iqzow6 = (Pqzow6 & Wqzow6);
assign Wqzow6 = (Drzow6 & Krzow6);
assign Krzow6 = (~(Fkfpw6[17] & Dfqow6));
assign Drzow6 = (Rrzow6 & Yrzow6);
assign Yrzow6 = (~(vis_psp_o[15] & Yfqow6));
assign Rrzow6 = (~(vis_msp_o[15] & Fgqow6));
assign Pqzow6 = (Fszow6 & Mszow6);
assign Mszow6 = (~(vis_r14_o[17] & Ahqow6));
assign Fszow6 = (~(vis_r12_o[17] & Hhqow6));
assign Bqzow6 = (Tszow6 & Atzow6);
assign Atzow6 = (Htzow6 & Otzow6);
assign Otzow6 = (~(vis_r9_o[17] & Qiqow6));
assign Htzow6 = (Vtzow6 & Cuzow6);
assign Cuzow6 = (~(vis_r11_o[17] & Ljqow6));
assign Vtzow6 = (~(vis_r10_o[17] & Sjqow6));
assign Tszow6 = (J10iu6 & Juzow6);
assign Juzow6 = (~(vis_r8_o[17] & Gkqow6));
assign J10iu6 = (Quzow6 & Xuzow6);
assign Xuzow6 = (Evzow6 & Lvzow6);
assign Lvzow6 = (Svzow6 & Zvzow6);
assign Zvzow6 = (~(vis_r2_o[17] & Dmqow6));
assign Svzow6 = (~(vis_r6_o[17] & Kmqow6));
assign Evzow6 = (Gwzow6 & Nwzow6);
assign Nwzow6 = (~(vis_r5_o[17] & Fnqow6));
assign Gwzow6 = (~(vis_r4_o[17] & Mnqow6));
assign Quzow6 = (Uwzow6 & Bxzow6);
assign Bxzow6 = (Ixzow6 & Pxzow6);
assign Pxzow6 = (~(vis_r1_o[17] & Voqow6));
assign Ixzow6 = (~(vis_r0_o[17] & Cpqow6));
assign Uwzow6 = (Wxzow6 & Dyzow6);
assign Dyzow6 = (~(vis_r3_o[17] & Xpqow6));
assign Wxzow6 = (~(vis_r7_o[17] & Eqqow6));
assign Gdqow6 = (Sevow6 & X71iu6);
assign Npzow6 = (~(G64iu6 & R0nhu6));
assign G64iu6 = (Shhpw6[17] & Iqzhu6);
assign HWDATA[15] = (~(Kyzow6 & Ryzow6));
assign Ryzow6 = (~(Yyzow6 & W89ju6));
assign W89ju6 = (~(Fzzow6 & Mzzow6));
assign Mzzow6 = (Tzzow6 & A00pw6);
assign A00pw6 = (H00pw6 & O00pw6);
assign O00pw6 = (~(Fkfpw6[15] & Dfqow6));
assign H00pw6 = (V00pw6 & C10pw6);
assign C10pw6 = (~(vis_psp_o[13] & Yfqow6));
assign V00pw6 = (~(vis_msp_o[13] & Fgqow6));
assign Tzzow6 = (J10pw6 & Q10pw6);
assign Q10pw6 = (~(vis_r14_o[15] & Ahqow6));
assign J10pw6 = (~(vis_r12_o[15] & Hhqow6));
assign Fzzow6 = (X10pw6 & E20pw6);
assign E20pw6 = (L20pw6 & S20pw6);
assign S20pw6 = (~(vis_r9_o[15] & Qiqow6));
assign L20pw6 = (Z20pw6 & G30pw6);
assign G30pw6 = (~(vis_r11_o[15] & Ljqow6));
assign Z20pw6 = (~(vis_r10_o[15] & Sjqow6));
assign X10pw6 = (X10iu6 & N30pw6);
assign N30pw6 = (~(vis_r8_o[15] & Gkqow6));
assign X10iu6 = (U30pw6 & B40pw6);
assign B40pw6 = (I40pw6 & P40pw6);
assign P40pw6 = (W40pw6 & D50pw6);
assign D50pw6 = (~(vis_r2_o[15] & Dmqow6));
assign W40pw6 = (~(vis_r6_o[15] & Kmqow6));
assign I40pw6 = (K50pw6 & R50pw6);
assign R50pw6 = (~(vis_r5_o[15] & Fnqow6));
assign K50pw6 = (~(vis_r4_o[15] & Mnqow6));
assign U30pw6 = (Y50pw6 & F60pw6);
assign F60pw6 = (M60pw6 & T60pw6);
assign T60pw6 = (~(vis_r1_o[15] & Voqow6));
assign M60pw6 = (~(vis_r0_o[15] & Cpqow6));
assign Y50pw6 = (A70pw6 & H70pw6);
assign H70pw6 = (~(vis_r3_o[15] & Xpqow6));
assign A70pw6 = (~(vis_r7_o[15] & Eqqow6));
assign Kyzow6 = (O70pw6 & Oqvow6);
assign Oqvow6 = (~(Udxow6 & Uo6ju6));
assign Uo6ju6 = (~(V70pw6 & C80pw6));
assign C80pw6 = (J80pw6 & Q80pw6);
assign Q80pw6 = (X80pw6 & E90pw6);
assign E90pw6 = (~(Fkfpw6[7] & Dfqow6));
assign X80pw6 = (L90pw6 & S90pw6);
assign S90pw6 = (~(vis_psp_o[5] & Yfqow6));
assign L90pw6 = (~(vis_msp_o[5] & Fgqow6));
assign J80pw6 = (Z90pw6 & Ga0pw6);
assign Ga0pw6 = (~(vis_r14_o[7] & Ahqow6));
assign Z90pw6 = (~(vis_r12_o[7] & Hhqow6));
assign V70pw6 = (Na0pw6 & Ua0pw6);
assign Ua0pw6 = (Bb0pw6 & Ib0pw6);
assign Ib0pw6 = (~(vis_r9_o[7] & Qiqow6));
assign Bb0pw6 = (Pb0pw6 & Wb0pw6);
assign Wb0pw6 = (~(vis_r11_o[7] & Ljqow6));
assign Pb0pw6 = (~(vis_r10_o[7] & Sjqow6));
assign Na0pw6 = (Svzhu6 & Dc0pw6);
assign Dc0pw6 = (~(vis_r8_o[7] & Gkqow6));
assign Svzhu6 = (Kc0pw6 & Rc0pw6);
assign Rc0pw6 = (Yc0pw6 & Fd0pw6);
assign Fd0pw6 = (Md0pw6 & Td0pw6);
assign Td0pw6 = (~(vis_r0_o[7] & Cpqow6));
assign Md0pw6 = (~(vis_r2_o[7] & Dmqow6));
assign Yc0pw6 = (Ae0pw6 & He0pw6);
assign He0pw6 = (~(vis_r5_o[7] & Fnqow6));
assign Ae0pw6 = (~(vis_r4_o[7] & Mnqow6));
assign Kc0pw6 = (Oe0pw6 & Ve0pw6);
assign Ve0pw6 = (Cf0pw6 & Jf0pw6);
assign Jf0pw6 = (~(vis_r7_o[7] & Eqqow6));
assign Cf0pw6 = (~(vis_r3_o[7] & Xpqow6));
assign Oe0pw6 = (Qf0pw6 & Xf0pw6);
assign Xf0pw6 = (~(vis_r1_o[7] & Voqow6));
assign Qf0pw6 = (~(vis_r6_o[7] & Kmqow6));
assign O70pw6 = (~(S54iu6 & R0nhu6));
assign S54iu6 = (Shhpw6[15] & Iqzhu6);
assign HWDATA[14] = (~(Eg0pw6 & Lg0pw6));
assign Lg0pw6 = (~(Yyzow6 & T39ju6));
assign T39ju6 = (~(Sg0pw6 & Zg0pw6));
assign Zg0pw6 = (Gh0pw6 & Nh0pw6);
assign Nh0pw6 = (Uh0pw6 & Bi0pw6);
assign Bi0pw6 = (~(vis_r11_o[14] & Ljqow6));
assign Uh0pw6 = (Ii0pw6 & Pi0pw6);
assign Pi0pw6 = (~(vis_r9_o[14] & Qiqow6));
assign Ii0pw6 = (~(Fkfpw6[14] & Dfqow6));
assign Gh0pw6 = (Wi0pw6 & Dj0pw6);
assign Dj0pw6 = (~(vis_r10_o[14] & Sjqow6));
assign Wi0pw6 = (~(vis_psp_o[12] & Yfqow6));
assign Sg0pw6 = (Kj0pw6 & Rj0pw6);
assign Rj0pw6 = (Yj0pw6 & Fk0pw6);
assign Fk0pw6 = (~(vis_r12_o[14] & Hhqow6));
assign Yj0pw6 = (Mk0pw6 & Tk0pw6);
assign Tk0pw6 = (~(vis_msp_o[12] & Fgqow6));
assign Mk0pw6 = (~(vis_r14_o[14] & Ahqow6));
assign Kj0pw6 = (E20iu6 & Al0pw6);
assign Al0pw6 = (~(vis_r8_o[14] & Gkqow6));
assign E20iu6 = (Hl0pw6 & Ol0pw6);
assign Ol0pw6 = (Vl0pw6 & Cm0pw6);
assign Cm0pw6 = (Jm0pw6 & Qm0pw6);
assign Qm0pw6 = (~(vis_r2_o[14] & Dmqow6));
assign Jm0pw6 = (~(vis_r6_o[14] & Kmqow6));
assign Vl0pw6 = (Xm0pw6 & En0pw6);
assign En0pw6 = (~(vis_r5_o[14] & Fnqow6));
assign Xm0pw6 = (~(vis_r4_o[14] & Mnqow6));
assign Hl0pw6 = (Ln0pw6 & Sn0pw6);
assign Sn0pw6 = (Zn0pw6 & Go0pw6);
assign Go0pw6 = (~(vis_r1_o[14] & Voqow6));
assign Zn0pw6 = (~(vis_r0_o[14] & Cpqow6));
assign Ln0pw6 = (No0pw6 & Uo0pw6);
assign Uo0pw6 = (~(vis_r3_o[14] & Xpqow6));
assign No0pw6 = (~(vis_r7_o[14] & Eqqow6));
assign Eg0pw6 = (Bp0pw6 & N0wow6);
assign N0wow6 = (~(Udxow6 & Kj6ju6));
assign Kj6ju6 = (~(Ip0pw6 & Pp0pw6));
assign Pp0pw6 = (Wp0pw6 & Dq0pw6);
assign Dq0pw6 = (Kq0pw6 & Rq0pw6);
assign Rq0pw6 = (~(Fkfpw6[6] & Dfqow6));
assign Kq0pw6 = (Yq0pw6 & Fr0pw6);
assign Fr0pw6 = (~(vis_psp_o[4] & Yfqow6));
assign Yq0pw6 = (~(vis_msp_o[4] & Fgqow6));
assign Wp0pw6 = (Mr0pw6 & Tr0pw6);
assign Tr0pw6 = (~(vis_r14_o[6] & Ahqow6));
assign Mr0pw6 = (~(vis_r12_o[6] & Hhqow6));
assign Ip0pw6 = (As0pw6 & Hs0pw6);
assign Hs0pw6 = (Os0pw6 & Vs0pw6);
assign Vs0pw6 = (~(vis_r9_o[6] & Qiqow6));
assign Os0pw6 = (Ct0pw6 & Jt0pw6);
assign Jt0pw6 = (~(vis_r11_o[6] & Ljqow6));
assign Ct0pw6 = (~(vis_r10_o[6] & Sjqow6));
assign As0pw6 = (Zvzhu6 & Qt0pw6);
assign Qt0pw6 = (~(vis_r8_o[6] & Gkqow6));
assign Zvzhu6 = (Xt0pw6 & Eu0pw6);
assign Eu0pw6 = (Lu0pw6 & Su0pw6);
assign Su0pw6 = (Zu0pw6 & Gv0pw6);
assign Gv0pw6 = (~(vis_r0_o[6] & Cpqow6));
assign Zu0pw6 = (~(vis_r2_o[6] & Dmqow6));
assign Lu0pw6 = (Nv0pw6 & Uv0pw6);
assign Uv0pw6 = (~(vis_r5_o[6] & Fnqow6));
assign Nv0pw6 = (~(vis_r4_o[6] & Mnqow6));
assign Xt0pw6 = (Bw0pw6 & Iw0pw6);
assign Iw0pw6 = (Pw0pw6 & Ww0pw6);
assign Ww0pw6 = (~(vis_r7_o[6] & Eqqow6));
assign Pw0pw6 = (~(vis_r3_o[6] & Xpqow6));
assign Bw0pw6 = (Dx0pw6 & Kx0pw6);
assign Kx0pw6 = (~(vis_r1_o[6] & Voqow6));
assign Dx0pw6 = (~(vis_r6_o[6] & Kmqow6));
assign Bp0pw6 = (~(L54iu6 & R0nhu6));
assign L54iu6 = (Shhpw6[14] & Iqzhu6);
assign HWDATA[13] = (~(Rx0pw6 & Yx0pw6));
assign Yx0pw6 = (~(Yyzow6 & Sz8ju6));
assign Sz8ju6 = (~(Fy0pw6 & My0pw6));
assign My0pw6 = (Ty0pw6 & Az0pw6);
assign Az0pw6 = (Hz0pw6 & Oz0pw6);
assign Oz0pw6 = (~(Fkfpw6[13] & Dfqow6));
assign Hz0pw6 = (Vz0pw6 & C01pw6);
assign C01pw6 = (~(vis_psp_o[11] & Yfqow6));
assign Vz0pw6 = (~(vis_msp_o[11] & Fgqow6));
assign Ty0pw6 = (J01pw6 & Q01pw6);
assign Q01pw6 = (~(vis_r14_o[13] & Ahqow6));
assign J01pw6 = (~(vis_r12_o[13] & Hhqow6));
assign Fy0pw6 = (X01pw6 & E11pw6);
assign E11pw6 = (L11pw6 & S11pw6);
assign S11pw6 = (~(vis_r9_o[13] & Qiqow6));
assign L11pw6 = (Z11pw6 & G21pw6);
assign G21pw6 = (~(vis_r11_o[13] & Ljqow6));
assign Z11pw6 = (~(vis_r10_o[13] & Sjqow6));
assign X01pw6 = (L20iu6 & N21pw6);
assign N21pw6 = (~(vis_r8_o[13] & Gkqow6));
assign L20iu6 = (U21pw6 & B31pw6);
assign B31pw6 = (I31pw6 & P31pw6);
assign P31pw6 = (W31pw6 & D41pw6);
assign D41pw6 = (~(vis_r2_o[13] & Dmqow6));
assign W31pw6 = (~(vis_r6_o[13] & Kmqow6));
assign I31pw6 = (K41pw6 & R41pw6);
assign R41pw6 = (~(vis_r5_o[13] & Fnqow6));
assign K41pw6 = (~(vis_r4_o[13] & Mnqow6));
assign U21pw6 = (Y41pw6 & F51pw6);
assign F51pw6 = (M51pw6 & T51pw6);
assign T51pw6 = (~(vis_r1_o[13] & Voqow6));
assign M51pw6 = (~(vis_r0_o[13] & Cpqow6));
assign Y41pw6 = (A61pw6 & H61pw6);
assign H61pw6 = (~(vis_r3_o[13] & Xpqow6));
assign A61pw6 = (~(vis_r7_o[13] & Eqqow6));
assign Rx0pw6 = (O61pw6 & Zqqow6);
assign Zqqow6 = (~(Udxow6 & Eg6ju6));
assign Eg6ju6 = (~(V61pw6 & C71pw6));
assign C71pw6 = (J71pw6 & Q71pw6);
assign Q71pw6 = (X71pw6 & E81pw6);
assign E81pw6 = (~(Fkfpw6[5] & Dfqow6));
assign X71pw6 = (L81pw6 & S81pw6);
assign S81pw6 = (~(vis_psp_o[3] & Yfqow6));
assign L81pw6 = (~(vis_msp_o[3] & Fgqow6));
assign J71pw6 = (Z81pw6 & G91pw6);
assign G91pw6 = (~(vis_r14_o[5] & Ahqow6));
assign Z81pw6 = (~(vis_r12_o[5] & Hhqow6));
assign V61pw6 = (N91pw6 & U91pw6);
assign U91pw6 = (Ba1pw6 & Ia1pw6);
assign Ia1pw6 = (~(vis_r9_o[5] & Qiqow6));
assign Ba1pw6 = (Pa1pw6 & Wa1pw6);
assign Wa1pw6 = (~(vis_r11_o[5] & Ljqow6));
assign Pa1pw6 = (~(vis_r10_o[5] & Sjqow6));
assign N91pw6 = (Gwzhu6 & Db1pw6);
assign Db1pw6 = (~(vis_r8_o[5] & Gkqow6));
assign Gwzhu6 = (Kb1pw6 & Rb1pw6);
assign Rb1pw6 = (Yb1pw6 & Fc1pw6);
assign Fc1pw6 = (Mc1pw6 & Tc1pw6);
assign Tc1pw6 = (~(vis_r0_o[5] & Cpqow6));
assign Mc1pw6 = (~(vis_r2_o[5] & Dmqow6));
assign Yb1pw6 = (Ad1pw6 & Hd1pw6);
assign Hd1pw6 = (~(vis_r5_o[5] & Fnqow6));
assign Ad1pw6 = (~(vis_r4_o[5] & Mnqow6));
assign Kb1pw6 = (Od1pw6 & Vd1pw6);
assign Vd1pw6 = (Ce1pw6 & Je1pw6);
assign Je1pw6 = (~(vis_r7_o[5] & Eqqow6));
assign Ce1pw6 = (~(vis_r3_o[5] & Xpqow6));
assign Od1pw6 = (Qe1pw6 & Xe1pw6);
assign Xe1pw6 = (~(vis_r1_o[5] & Voqow6));
assign Qe1pw6 = (~(vis_r6_o[5] & Kmqow6));
assign O61pw6 = (~(E54iu6 & R0nhu6));
assign E54iu6 = (Shhpw6[13] & Iqzhu6);
assign HWDATA[12] = (~(Ef1pw6 & Lf1pw6));
assign Lf1pw6 = (~(Yyzow6 & Rv8ju6));
assign Rv8ju6 = (~(Sf1pw6 & Zf1pw6));
assign Zf1pw6 = (Gg1pw6 & Ng1pw6);
assign Ng1pw6 = (Ug1pw6 & Bh1pw6);
assign Bh1pw6 = (~(vis_r11_o[12] & Ljqow6));
assign Ug1pw6 = (Ih1pw6 & Ph1pw6);
assign Ph1pw6 = (~(vis_r10_o[12] & Sjqow6));
assign Ih1pw6 = (~(vis_r9_o[12] & Qiqow6));
assign Gg1pw6 = (Wh1pw6 & Di1pw6);
assign Di1pw6 = (~(Fkfpw6[12] & Dfqow6));
assign Wh1pw6 = (~(vis_r12_o[12] & Hhqow6));
assign Sf1pw6 = (Ki1pw6 & Ri1pw6);
assign Ri1pw6 = (Yi1pw6 & Fj1pw6);
assign Fj1pw6 = (~(vis_r14_o[12] & Ahqow6));
assign Yi1pw6 = (Mj1pw6 & Tj1pw6);
assign Tj1pw6 = (~(vis_psp_o[10] & Yfqow6));
assign Mj1pw6 = (~(vis_r8_o[12] & Gkqow6));
assign Ki1pw6 = (S20iu6 & Ak1pw6);
assign Ak1pw6 = (~(vis_msp_o[10] & Fgqow6));
assign S20iu6 = (Hk1pw6 & Ok1pw6);
assign Ok1pw6 = (Vk1pw6 & Cl1pw6);
assign Cl1pw6 = (Jl1pw6 & Ql1pw6);
assign Ql1pw6 = (~(vis_r0_o[12] & Cpqow6));
assign Jl1pw6 = (~(vis_r2_o[12] & Dmqow6));
assign Vk1pw6 = (Xl1pw6 & Em1pw6);
assign Em1pw6 = (~(vis_r5_o[12] & Fnqow6));
assign Xl1pw6 = (~(vis_r4_o[12] & Mnqow6));
assign Hk1pw6 = (Lm1pw6 & Sm1pw6);
assign Sm1pw6 = (Zm1pw6 & Gn1pw6);
assign Gn1pw6 = (~(vis_r7_o[12] & Eqqow6));
assign Zm1pw6 = (~(vis_r3_o[12] & Xpqow6));
assign Lm1pw6 = (Nn1pw6 & Un1pw6);
assign Un1pw6 = (~(vis_r1_o[12] & Voqow6));
assign Nn1pw6 = (~(vis_r6_o[12] & Kmqow6));
assign Ef1pw6 = (Bo1pw6 & Abwow6);
assign Abwow6 = (~(Udxow6 & Zw4ju6));
assign Zw4ju6 = (~(Io1pw6 & Po1pw6));
assign Po1pw6 = (Wo1pw6 & Dp1pw6);
assign Dp1pw6 = (Kp1pw6 & Rp1pw6);
assign Rp1pw6 = (~(Fkfpw6[4] & Dfqow6));
assign Kp1pw6 = (Yp1pw6 & Fq1pw6);
assign Fq1pw6 = (~(vis_psp_o[2] & Yfqow6));
assign Yp1pw6 = (~(vis_msp_o[2] & Fgqow6));
assign Wo1pw6 = (Mq1pw6 & Tq1pw6);
assign Tq1pw6 = (~(vis_r14_o[4] & Ahqow6));
assign Mq1pw6 = (~(vis_r12_o[4] & Hhqow6));
assign Io1pw6 = (Ar1pw6 & Hr1pw6);
assign Hr1pw6 = (Or1pw6 & Vr1pw6);
assign Vr1pw6 = (~(vis_r9_o[4] & Qiqow6));
assign Or1pw6 = (Cs1pw6 & Js1pw6);
assign Js1pw6 = (~(vis_r11_o[4] & Ljqow6));
assign Cs1pw6 = (~(vis_r10_o[4] & Sjqow6));
assign Ar1pw6 = (Nwzhu6 & Qs1pw6);
assign Qs1pw6 = (~(vis_r8_o[4] & Gkqow6));
assign Nwzhu6 = (Xs1pw6 & Et1pw6);
assign Et1pw6 = (Lt1pw6 & St1pw6);
assign St1pw6 = (Zt1pw6 & Gu1pw6);
assign Gu1pw6 = (~(vis_r0_o[4] & Cpqow6));
assign Zt1pw6 = (~(vis_r2_o[4] & Dmqow6));
assign Lt1pw6 = (Nu1pw6 & Uu1pw6);
assign Uu1pw6 = (~(vis_r5_o[4] & Fnqow6));
assign Nu1pw6 = (~(vis_r4_o[4] & Mnqow6));
assign Xs1pw6 = (Bv1pw6 & Iv1pw6);
assign Iv1pw6 = (Pv1pw6 & Wv1pw6);
assign Wv1pw6 = (~(vis_r7_o[4] & Eqqow6));
assign Pv1pw6 = (~(vis_r3_o[4] & Xpqow6));
assign Bv1pw6 = (Dw1pw6 & Kw1pw6);
assign Kw1pw6 = (~(vis_r1_o[4] & Voqow6));
assign Dw1pw6 = (~(vis_r6_o[4] & Kmqow6));
assign Bo1pw6 = (~(X44iu6 & R0nhu6));
assign X44iu6 = (Shhpw6[12] & Iqzhu6);
assign HWDATA[11] = (~(Rw1pw6 & Yw1pw6));
assign Yw1pw6 = (~(Yyzow6 & In8ju6));
assign In8ju6 = (~(Fx1pw6 & Mx1pw6));
assign Mx1pw6 = (Tx1pw6 & Ay1pw6);
assign Ay1pw6 = (Hy1pw6 & Oy1pw6);
assign Oy1pw6 = (~(vis_r11_o[11] & Ljqow6));
assign Hy1pw6 = (Vy1pw6 & Cz1pw6);
assign Cz1pw6 = (~(vis_r9_o[11] & Qiqow6));
assign Vy1pw6 = (~(Fkfpw6[11] & Dfqow6));
assign Tx1pw6 = (Jz1pw6 & Qz1pw6);
assign Qz1pw6 = (~(vis_r10_o[11] & Sjqow6));
assign Jz1pw6 = (~(vis_psp_o[9] & Yfqow6));
assign Fx1pw6 = (Xz1pw6 & E02pw6);
assign E02pw6 = (L02pw6 & S02pw6);
assign S02pw6 = (~(vis_r12_o[11] & Hhqow6));
assign L02pw6 = (Z02pw6 & G12pw6);
assign G12pw6 = (~(vis_msp_o[9] & Fgqow6));
assign Z02pw6 = (~(vis_r14_o[11] & Ahqow6));
assign Xz1pw6 = (Z20iu6 & N12pw6);
assign N12pw6 = (~(vis_r8_o[11] & Gkqow6));
assign Z20iu6 = (U12pw6 & B22pw6);
assign B22pw6 = (I22pw6 & P22pw6);
assign P22pw6 = (W22pw6 & D32pw6);
assign D32pw6 = (~(vis_r2_o[11] & Dmqow6));
assign W22pw6 = (~(vis_r6_o[11] & Kmqow6));
assign I22pw6 = (K32pw6 & R32pw6);
assign R32pw6 = (~(vis_r5_o[11] & Fnqow6));
assign K32pw6 = (~(vis_r4_o[11] & Mnqow6));
assign U12pw6 = (Y32pw6 & F42pw6);
assign F42pw6 = (M42pw6 & T42pw6);
assign T42pw6 = (~(vis_r1_o[11] & Voqow6));
assign M42pw6 = (~(vis_r0_o[11] & Cpqow6));
assign Y32pw6 = (A52pw6 & H52pw6);
assign H52pw6 = (~(vis_r3_o[11] & Xpqow6));
assign A52pw6 = (~(vis_r7_o[11] & Eqqow6));
assign Rw1pw6 = (O52pw6 & Zkwow6);
assign Zkwow6 = (~(Udxow6 & G36ju6));
assign G36ju6 = (~(V52pw6 & C62pw6));
assign C62pw6 = (J62pw6 & Q62pw6);
assign Q62pw6 = (X62pw6 & E72pw6);
assign E72pw6 = (~(Fkfpw6[3] & Dfqow6));
assign X62pw6 = (L72pw6 & S72pw6);
assign S72pw6 = (~(vis_psp_o[1] & Yfqow6));
assign L72pw6 = (~(vis_msp_o[1] & Fgqow6));
assign J62pw6 = (Z72pw6 & G82pw6);
assign G82pw6 = (~(vis_r14_o[3] & Ahqow6));
assign Z72pw6 = (~(vis_r12_o[3] & Hhqow6));
assign V52pw6 = (N82pw6 & U82pw6);
assign U82pw6 = (B92pw6 & I92pw6);
assign I92pw6 = (~(vis_r9_o[3] & Qiqow6));
assign B92pw6 = (P92pw6 & W92pw6);
assign W92pw6 = (~(vis_r11_o[3] & Ljqow6));
assign P92pw6 = (~(vis_r10_o[3] & Sjqow6));
assign N82pw6 = (Uwzhu6 & Da2pw6);
assign Da2pw6 = (~(vis_r8_o[3] & Gkqow6));
assign Uwzhu6 = (Ka2pw6 & Ra2pw6);
assign Ra2pw6 = (Ya2pw6 & Fb2pw6);
assign Fb2pw6 = (Mb2pw6 & Tb2pw6);
assign Tb2pw6 = (~(vis_r0_o[3] & Cpqow6));
assign Mb2pw6 = (~(vis_r2_o[3] & Dmqow6));
assign Ya2pw6 = (Ac2pw6 & Hc2pw6);
assign Hc2pw6 = (~(vis_r5_o[3] & Fnqow6));
assign Ac2pw6 = (~(vis_r4_o[3] & Mnqow6));
assign Ka2pw6 = (Oc2pw6 & Vc2pw6);
assign Vc2pw6 = (Cd2pw6 & Jd2pw6);
assign Jd2pw6 = (~(vis_r7_o[3] & Eqqow6));
assign Cd2pw6 = (~(vis_r3_o[3] & Xpqow6));
assign Oc2pw6 = (Qd2pw6 & Xd2pw6);
assign Xd2pw6 = (~(vis_r1_o[3] & Voqow6));
assign Qd2pw6 = (~(vis_r6_o[3] & Kmqow6));
assign O52pw6 = (~(Q44iu6 & R0nhu6));
assign Q44iu6 = (Shhpw6[11] & Iqzhu6);
assign HWDATA[10] = (~(Ee2pw6 & Le2pw6));
assign Le2pw6 = (Vcvow6 | Ka8ju6);
assign Ka8ju6 = (Se2pw6 & Ze2pw6);
assign Ze2pw6 = (Gf2pw6 & Nf2pw6);
assign Nf2pw6 = (Uf2pw6 & Bg2pw6);
assign Bg2pw6 = (~(vis_r11_o[10] & Ljqow6));
assign Uf2pw6 = (Ig2pw6 & Pg2pw6);
assign Pg2pw6 = (~(vis_r9_o[10] & Qiqow6));
assign Ig2pw6 = (~(Fkfpw6[10] & Dfqow6));
assign Gf2pw6 = (Wg2pw6 & Dh2pw6);
assign Dh2pw6 = (~(vis_r10_o[10] & Sjqow6));
assign Wg2pw6 = (~(vis_psp_o[8] & Yfqow6));
assign Se2pw6 = (Kh2pw6 & Rh2pw6);
assign Rh2pw6 = (Yh2pw6 & Fi2pw6);
assign Fi2pw6 = (~(vis_r12_o[10] & Hhqow6));
assign Yh2pw6 = (Mi2pw6 & Ti2pw6);
assign Ti2pw6 = (~(vis_msp_o[8] & Fgqow6));
assign Mi2pw6 = (~(vis_r14_o[10] & Ahqow6));
assign Kh2pw6 = (G30iu6 & Aj2pw6);
assign Aj2pw6 = (~(vis_r8_o[10] & Gkqow6));
assign G30iu6 = (Hj2pw6 & Oj2pw6);
assign Oj2pw6 = (Vj2pw6 & Ck2pw6);
assign Ck2pw6 = (Jk2pw6 & Qk2pw6);
assign Qk2pw6 = (~(vis_r2_o[10] & Dmqow6));
assign Jk2pw6 = (~(vis_r6_o[10] & Kmqow6));
assign Vj2pw6 = (Xk2pw6 & El2pw6);
assign El2pw6 = (~(vis_r5_o[10] & Fnqow6));
assign Xk2pw6 = (~(vis_r4_o[10] & Mnqow6));
assign Hj2pw6 = (Ll2pw6 & Sl2pw6);
assign Sl2pw6 = (Zl2pw6 & Gm2pw6);
assign Gm2pw6 = (~(vis_r1_o[10] & Voqow6));
assign Zl2pw6 = (~(vis_r0_o[10] & Cpqow6));
assign Ll2pw6 = (Nm2pw6 & Um2pw6);
assign Um2pw6 = (~(vis_r3_o[10] & Xpqow6));
assign Nm2pw6 = (~(vis_r7_o[10] & Eqqow6));
assign Vcvow6 = (!Yyzow6);
assign Yyzow6 = (Qaxiu6 & Bn2pw6);
assign Bn2pw6 = (~(J71iu6 & L3ehu6));
assign Ee2pw6 = (In2pw6 & Fvwow6);
assign Fvwow6 = (~(Udxow6 & Ot5ju6));
assign Ot5ju6 = (~(Pn2pw6 & Wn2pw6));
assign Wn2pw6 = (Do2pw6 & Ko2pw6);
assign Ko2pw6 = (Ro2pw6 & Yo2pw6);
assign Yo2pw6 = (~(Fkfpw6[2] & Dfqow6));
assign Ro2pw6 = (Fp2pw6 & Mp2pw6);
assign Mp2pw6 = (~(vis_psp_o[0] & Yfqow6));
assign Yfqow6 = (Tp2pw6 & Vrfhu6);
assign Tp2pw6 = (Aq2pw6 & Hq2pw6);
assign Fp2pw6 = (~(vis_msp_o[0] & Fgqow6));
assign Fgqow6 = (Oq2pw6 & Aq2pw6);
assign Oq2pw6 = (Hq2pw6 & Vq2pw6);
assign Do2pw6 = (Cr2pw6 & Jr2pw6);
assign Jr2pw6 = (~(vis_r14_o[2] & Ahqow6));
assign Cr2pw6 = (~(vis_r12_o[2] & Hhqow6));
assign Pn2pw6 = (Qr2pw6 & Xr2pw6);
assign Xr2pw6 = (Es2pw6 & Ls2pw6);
assign Ls2pw6 = (~(vis_r9_o[2] & Qiqow6));
assign Es2pw6 = (Ss2pw6 & Zs2pw6);
assign Zs2pw6 = (~(vis_r11_o[2] & Ljqow6));
assign Ss2pw6 = (~(vis_r10_o[2] & Sjqow6));
assign Qr2pw6 = (Pxzhu6 & Gt2pw6);
assign Gt2pw6 = (~(vis_r8_o[2] & Gkqow6));
assign Pxzhu6 = (Nt2pw6 & Ut2pw6);
assign Ut2pw6 = (Bu2pw6 & Iu2pw6);
assign Iu2pw6 = (Pu2pw6 & Wu2pw6);
assign Wu2pw6 = (~(vis_r0_o[2] & Cpqow6));
assign Pu2pw6 = (~(vis_r2_o[2] & Dmqow6));
assign Bu2pw6 = (Dv2pw6 & Kv2pw6);
assign Kv2pw6 = (~(vis_r5_o[2] & Fnqow6));
assign Dv2pw6 = (~(vis_r4_o[2] & Mnqow6));
assign Nt2pw6 = (Rv2pw6 & Yv2pw6);
assign Yv2pw6 = (Fw2pw6 & Mw2pw6);
assign Mw2pw6 = (~(vis_r7_o[2] & Eqqow6));
assign Fw2pw6 = (~(vis_r3_o[2] & Xpqow6));
assign Rv2pw6 = (Tw2pw6 & Ax2pw6);
assign Ax2pw6 = (~(vis_r1_o[2] & Voqow6));
assign Tw2pw6 = (~(vis_r6_o[2] & Kmqow6));
assign Udxow6 = (J71iu6 & Sevow6);
assign In2pw6 = (~(J44iu6 & R0nhu6));
assign J44iu6 = (Shhpw6[10] & Iqzhu6);
assign HWDATA[0] = (~(Hx2pw6 & Ox2pw6));
assign Ox2pw6 = (~(Sevow6 & L35ju6));
assign L35ju6 = (~(Vx2pw6 & Cy2pw6));
assign Cy2pw6 = (Jy2pw6 & Qy2pw6);
assign Qy2pw6 = (Xy2pw6 & Ez2pw6);
assign Ez2pw6 = (~(Fkfpw6[0] & Dfqow6));
assign Dfqow6 = (Lz2pw6 & Aq2pw6);
assign Xy2pw6 = (~(vis_r14_o[0] & Ahqow6));
assign Ahqow6 = (Sz2pw6 & Aq2pw6);
assign Jy2pw6 = (Zz2pw6 & G03pw6);
assign G03pw6 = (~(vis_r12_o[0] & Hhqow6));
assign Hhqow6 = (Aq2pw6 & N03pw6);
assign Aq2pw6 = (~(Ntniu6 | Roniu6));
assign Zz2pw6 = (~(vis_r11_o[0] & Ljqow6));
assign Ljqow6 = (Lz2pw6 & U03pw6);
assign Lz2pw6 = (~(Qrniu6 | Ivuow6));
assign Vx2pw6 = (B13pw6 & I13pw6);
assign I13pw6 = (P13pw6 & W13pw6);
assign W13pw6 = (~(vis_r10_o[0] & Sjqow6));
assign Sjqow6 = (Sz2pw6 & U03pw6);
assign Sz2pw6 = (~(Ivuow6 | X3fpw6[0]));
assign P13pw6 = (~(vis_r9_o[0] & Qiqow6));
assign Qiqow6 = (U03pw6 & Hq2pw6);
assign B13pw6 = (N30iu6 & D23pw6);
assign D23pw6 = (~(vis_r8_o[0] & Gkqow6));
assign Gkqow6 = (U03pw6 & N03pw6);
assign U03pw6 = (~(Ntniu6 | X3fpw6[2]));
assign Ntniu6 = (!X3fpw6[3]);
assign N30iu6 = (K23pw6 & R23pw6);
assign R23pw6 = (Y23pw6 & F33pw6);
assign F33pw6 = (M33pw6 & T33pw6);
assign T33pw6 = (~(vis_r0_o[0] & Cpqow6));
assign Cpqow6 = (A43pw6 & N03pw6);
assign M33pw6 = (~(vis_r2_o[0] & Dmqow6));
assign Dmqow6 = (H43pw6 & O43pw6);
assign H43pw6 = (~(X3fpw6[0] | X3fpw6[2]));
assign Y23pw6 = (V43pw6 & C53pw6);
assign C53pw6 = (~(vis_r5_o[0] & Fnqow6));
assign Fnqow6 = (J53pw6 & Hq2pw6);
assign V43pw6 = (~(vis_r4_o[0] & Mnqow6));
assign Mnqow6 = (J53pw6 & N03pw6);
assign N03pw6 = (~(X3fpw6[0] | X3fpw6[1]));
assign J53pw6 = (~(Roniu6 | X3fpw6[3]));
assign K23pw6 = (Q53pw6 & X53pw6);
assign X53pw6 = (E63pw6 & L63pw6);
assign L63pw6 = (~(vis_r7_o[0] & Eqqow6));
assign Eqqow6 = (S63pw6 & X3fpw6[0]);
assign S63pw6 = (X3fpw6[2] & O43pw6);
assign E63pw6 = (~(vis_r3_o[0] & Xpqow6));
assign Xpqow6 = (Z63pw6 & X3fpw6[0]);
assign Z63pw6 = (O43pw6 & Roniu6);
assign Roniu6 = (!X3fpw6[2]);
assign Q53pw6 = (G73pw6 & N73pw6);
assign N73pw6 = (~(vis_r1_o[0] & Voqow6));
assign Voqow6 = (A43pw6 & Hq2pw6);
assign Hq2pw6 = (~(Qrniu6 | X3fpw6[1]));
assign A43pw6 = (~(X3fpw6[2] | X3fpw6[3]));
assign G73pw6 = (~(vis_r6_o[0] & Kmqow6));
assign Kmqow6 = (U73pw6 & X3fpw6[2]);
assign U73pw6 = (O43pw6 & Qrniu6);
assign Qrniu6 = (!X3fpw6[0]);
assign O43pw6 = (~(Ivuow6 | X3fpw6[3]));
assign Ivuow6 = (!X3fpw6[1]);
assign Sevow6 = (L3ehu6 & Qaxiu6);
assign Qaxiu6 = (!R0nhu6);
assign Hx2pw6 = (~(T24iu6 & R0nhu6));
assign T24iu6 = (Shhpw6[0] & Iqzhu6);
assign HTRANS[1] = (~(B83pw6 & I83pw6));
assign I83pw6 = (~(Xg6iu6 & Kzciu6));
assign Kzciu6 = (~(P83pw6 & W83pw6));
assign W83pw6 = (~(D93pw6 | Jshpw6[28]));
assign D93pw6 = (!Jshpw6[31]);
assign P83pw6 = (Jshpw6[30] & Jshpw6[29]);
assign B83pw6 = (W7cow6 ? I7cow6 : K93pw6);
assign W7cow6 = (Ympiu6 & L18iu6);
assign I7cow6 = (Dx0iu6 ? Ef1iu6 : Rx0iu6);
assign K93pw6 = (~(R93pw6 & S18iu6));
assign R93pw6 = (Y93pw6 & Z18iu6);
assign Z18iu6 = (~(Fa3pw6 & Ma3pw6));
assign Ma3pw6 = (~(Ta3pw6 & Ab3pw6));
assign Ab3pw6 = (~(Iiliu6 & Hb3pw6));
assign Hb3pw6 = (X71iu6 | Ympiu6);
assign Fa3pw6 = (~(J71iu6 & Ob3pw6));
assign Y93pw6 = (Pyciu6 | V0epw6);
assign Pyciu6 = (~(Vb3pw6 & Ef1iu6));
assign Vb3pw6 = (Rx0iu6 & Dx0iu6);
assign HSIZE[1] = (!Cc3pw6);
assign Cc3pw6 = (Xg6iu6 ? Qc3pw6 : Jc3pw6);
assign Qc3pw6 = (~(Aphpw6[2] | Wqzhu6));
assign Jc3pw6 = (Ob3pw6 & Xc3pw6);
assign Xc3pw6 = (Ed3pw6 | Sdaiu6);
assign HSIZE[0] = (~(Ld3pw6 & Sd3pw6));
assign Sd3pw6 = (~(Zd3pw6 & Ge3pw6));
assign Ge3pw6 = (~(Ympiu6 | Sdaiu6));
assign Zd3pw6 = (Mnxow6 & Ze9iu6);
assign Ld3pw6 = (~(Ne3pw6 & Aphpw6[1]));
assign HPROT[3] = (~(HPROT[2] & Ue3pw6));
assign Ue3pw6 = (~(HADDR[29] & Bf3pw6));
assign Bf3pw6 = (!HADDR[31]);
assign HADDR[31] = (Xg6iu6 ? Jshpw6[31] : Ef1iu6);
assign Ef1iu6 = (~(If3pw6 & Pf3pw6));
assign Pf3pw6 = (T2iiu6 | R65ju6);
assign R65ju6 = (Mm4ju6 ? Wf3pw6 : Wtoiu6);
assign Wf3pw6 = (Dg3pw6 & Kg3pw6);
assign Kg3pw6 = (Rg3pw6 & Yg3pw6);
assign Yg3pw6 = (Fh3pw6 & Mh3pw6);
assign Mh3pw6 = (~(Jo4ju6 & vis_r14_o[31]));
assign Fh3pw6 = (Th3pw6 & Ai3pw6);
assign Ai3pw6 = (~(Ep4ju6 & vis_psp_o[29]));
assign Th3pw6 = (~(Lp4ju6 & vis_msp_o[29]));
assign Rg3pw6 = (Hi3pw6 & Oi3pw6);
assign Oi3pw6 = (~(Gq4ju6 & vis_r12_o[31]));
assign Hi3pw6 = (~(Nq4ju6 & vis_r11_o[31]));
assign Dg3pw6 = (Vi3pw6 & Cj3pw6);
assign Cj3pw6 = (Jj3pw6 & Qj3pw6);
assign Qj3pw6 = (~(Wr4ju6 & vis_r10_o[31]));
assign Jj3pw6 = (~(Ds4ju6 & vis_r9_o[31]));
assign Vi3pw6 = (R50iu6 & Xj3pw6);
assign Xj3pw6 = (~(Rs4ju6 & vis_r8_o[31]));
assign R50iu6 = (Ek3pw6 & Lk3pw6);
assign Lk3pw6 = (Sk3pw6 & Zk3pw6);
assign Zk3pw6 = (Gl3pw6 & Nl3pw6);
assign Nl3pw6 = (~(V6now6 & vis_r2_o[31]));
assign Gl3pw6 = (~(C7now6 & vis_r6_o[31]));
assign Sk3pw6 = (Ul3pw6 & Bm3pw6);
assign Bm3pw6 = (~(X7now6 & vis_r5_o[31]));
assign Ul3pw6 = (~(E8now6 & vis_r4_o[31]));
assign Ek3pw6 = (Im3pw6 & Pm3pw6);
assign Pm3pw6 = (Wm3pw6 & Dn3pw6);
assign Dn3pw6 = (~(N9now6 & vis_r1_o[31]));
assign Wm3pw6 = (~(U9now6 & vis_r0_o[31]));
assign Im3pw6 = (Kn3pw6 & Rn3pw6);
assign Rn3pw6 = (~(Panow6 & vis_r3_o[31]));
assign Kn3pw6 = (~(Wanow6 & vis_r7_o[31]));
assign Wtoiu6 = (!Fkfpw6[31]);
assign If3pw6 = (Yn3pw6 & Fo3pw6);
assign Fo3pw6 = (~(Eafpw6[31] & A3iiu6));
assign Yn3pw6 = (~(N5fpw6[30] & Sdaiu6));
assign HPROT[2] = (HADDR[30] | HADDR[29]);
assign HPROT[0] = (~(L18iu6 & Ze9iu6));
assign L18iu6 = (Mo3pw6 & To3pw6);
assign To3pw6 = (Ap3pw6 & Hp3pw6);
assign Hp3pw6 = (Op3pw6 & Hq1ju6);
assign Hq1ju6 = (~(Vp3pw6 & Pthiu6));
assign Vp3pw6 = (Ls1ju6 & Y2oiu6);
assign Op3pw6 = (Cq3pw6 & Oq1ju6);
assign Ap3pw6 = (Jq3pw6 & Qq3pw6);
assign Qq3pw6 = (~(Xq3pw6 & Glaiu6));
assign Glaiu6 = (M2piu6 & Cyfpw6[5]);
assign M2piu6 = (Xzmiu6 & Y7ghu6);
assign Xq3pw6 = (~(Mmjiu6 | Ae0iu6));
assign Jq3pw6 = (Bgaow6 & Er3pw6);
assign Er3pw6 = (~(I82ju6 & Oiaiu6));
assign Bgaow6 = (~(Lr3pw6 & Whfiu6));
assign Lr3pw6 = (D6kiu6 & Sijiu6);
assign Mo3pw6 = (Sr3pw6 & Zr3pw6);
assign Zr3pw6 = (Gs3pw6 & Ns3pw6);
assign Ns3pw6 = (~(Qe8iu6 & Us3pw6));
assign Us3pw6 = (~(S62ju6 & Jc2ju6));
assign S62ju6 = (Mr0iu6 | Cyfpw6[4]);
assign Gs3pw6 = (Bt3pw6 & It3pw6);
assign It3pw6 = (~(Y0jiu6 & Zqaju6));
assign Zqaju6 = (Sijiu6 & Ii0iu6);
assign Bt3pw6 = (~(Pt3pw6 & O96ow6));
assign O96ow6 = (Cyfpw6[4] & Geaiu6);
assign Pt3pw6 = (~(R2aiu6 | Cyfpw6[6]));
assign Sr3pw6 = (Yavow6 & Rcziu6);
assign Yavow6 = (Wt3pw6 & Du3pw6);
assign Du3pw6 = (~(Ku3pw6 & Mo2ju6));
assign Mo2ju6 = (Nlaiu6 & Hs0iu6);
assign Ku3pw6 = (~(P1bow6 | Cyfpw6[4]));
assign Wt3pw6 = (~(Ru3pw6 & Apaiu6));
assign Ru3pw6 = (~(Lkaiu6 | Mr0iu6));
assign HALTED = (Pzwiu6 & Wofiu6);
assign HADDR[9] = (Xg6iu6 ? Jshpw6[9] : Tugpw6[7]);
assign Tugpw6[7] = (~(Yu3pw6 & Fv3pw6));
assign Fv3pw6 = (~(N5fpw6[8] & Sdaiu6));
assign Yu3pw6 = (Mv3pw6 & Tv3pw6);
assign Tv3pw6 = (~(B7iiu6 & He0iu6));
assign He0iu6 = (Cn5ju6 ? Fkfpw6[9] : Aw3pw6);
assign Aw3pw6 = (~(Hw3pw6 & Ow3pw6));
assign Ow3pw6 = (Vw3pw6 & Cx3pw6);
assign Cx3pw6 = (Jx3pw6 & Qx3pw6);
assign Qx3pw6 = (~(Jo4ju6 & vis_r14_o[9]));
assign Jx3pw6 = (Xx3pw6 & Ey3pw6);
assign Ey3pw6 = (~(Ep4ju6 & vis_psp_o[7]));
assign Xx3pw6 = (~(Lp4ju6 & vis_msp_o[7]));
assign Vw3pw6 = (Ly3pw6 & Sy3pw6);
assign Sy3pw6 = (~(Gq4ju6 & vis_r12_o[9]));
assign Ly3pw6 = (~(Nq4ju6 & vis_r11_o[9]));
assign Hw3pw6 = (Zy3pw6 & Gz3pw6);
assign Gz3pw6 = (Nz3pw6 & Uz3pw6);
assign Uz3pw6 = (~(Wr4ju6 & vis_r10_o[9]));
assign Nz3pw6 = (~(Ds4ju6 & vis_r9_o[9]));
assign Zy3pw6 = (U30iu6 & B04pw6);
assign B04pw6 = (~(Rs4ju6 & vis_r8_o[9]));
assign U30iu6 = (I04pw6 & P04pw6);
assign P04pw6 = (W04pw6 & D14pw6);
assign D14pw6 = (K14pw6 & R14pw6);
assign R14pw6 = (~(V6now6 & vis_r2_o[9]));
assign K14pw6 = (~(C7now6 & vis_r6_o[9]));
assign W04pw6 = (Y14pw6 & F24pw6);
assign F24pw6 = (~(X7now6 & vis_r5_o[9]));
assign Y14pw6 = (~(E8now6 & vis_r4_o[9]));
assign I04pw6 = (M24pw6 & T24pw6);
assign T24pw6 = (A34pw6 & H34pw6);
assign H34pw6 = (~(N9now6 & vis_r1_o[9]));
assign A34pw6 = (~(U9now6 & vis_r0_o[9]));
assign M24pw6 = (O34pw6 & V34pw6);
assign V34pw6 = (~(Panow6 & vis_r3_o[9]));
assign O34pw6 = (~(Wanow6 & vis_r7_o[9]));
assign Mv3pw6 = (~(Eafpw6[9] & A3iiu6));
assign HADDR[6] = (Xg6iu6 ? Jshpw6[6] : Tugpw6[4]);
assign Tugpw6[4] = (~(C44pw6 & J44pw6));
assign J44pw6 = (~(N5fpw6[5] & Sdaiu6));
assign C44pw6 = (Q44pw6 & X44pw6);
assign X44pw6 = (~(B7iiu6 & Qf0iu6));
assign Qf0iu6 = (Cn5ju6 ? Fkfpw6[6] : E54pw6);
assign E54pw6 = (~(L54pw6 & S54pw6));
assign S54pw6 = (Z54pw6 & G64pw6);
assign G64pw6 = (N64pw6 & U64pw6);
assign U64pw6 = (~(Jo4ju6 & vis_r14_o[6]));
assign N64pw6 = (B74pw6 & I74pw6);
assign I74pw6 = (~(Ep4ju6 & vis_psp_o[4]));
assign B74pw6 = (~(Lp4ju6 & vis_msp_o[4]));
assign Z54pw6 = (P74pw6 & W74pw6);
assign W74pw6 = (~(Gq4ju6 & vis_r12_o[6]));
assign P74pw6 = (~(Nq4ju6 & vis_r11_o[6]));
assign L54pw6 = (D84pw6 & K84pw6);
assign K84pw6 = (R84pw6 & Y84pw6);
assign Y84pw6 = (~(Wr4ju6 & vis_r10_o[6]));
assign R84pw6 = (~(Ds4ju6 & vis_r9_o[6]));
assign D84pw6 = (P40iu6 & F94pw6);
assign F94pw6 = (~(Rs4ju6 & vis_r8_o[6]));
assign P40iu6 = (M94pw6 & T94pw6);
assign T94pw6 = (Aa4pw6 & Ha4pw6);
assign Ha4pw6 = (Oa4pw6 & Va4pw6);
assign Va4pw6 = (~(V6now6 & vis_r2_o[6]));
assign Oa4pw6 = (~(C7now6 & vis_r6_o[6]));
assign Aa4pw6 = (Cb4pw6 & Jb4pw6);
assign Jb4pw6 = (~(X7now6 & vis_r5_o[6]));
assign Cb4pw6 = (~(E8now6 & vis_r4_o[6]));
assign M94pw6 = (Qb4pw6 & Xb4pw6);
assign Xb4pw6 = (Ec4pw6 & Lc4pw6);
assign Lc4pw6 = (~(N9now6 & vis_r1_o[6]));
assign Ec4pw6 = (~(U9now6 & vis_r0_o[6]));
assign Qb4pw6 = (Sc4pw6 & Zc4pw6);
assign Zc4pw6 = (~(Panow6 & vis_r3_o[6]));
assign Sc4pw6 = (~(Wanow6 & vis_r7_o[6]));
assign Q44pw6 = (~(Eafpw6[6] & A3iiu6));
assign HADDR[30] = (Ze9iu6 ? Rx0iu6 : Jshpw6[30]);
assign Rx0iu6 = (~(Gd4pw6 & Nd4pw6));
assign Nd4pw6 = (T2iiu6 | Sg0iu6);
assign Sg0iu6 = (Mm4ju6 ? Ud4pw6 : Galiu6);
assign Ud4pw6 = (Be4pw6 & Ie4pw6);
assign Ie4pw6 = (Pe4pw6 & We4pw6);
assign We4pw6 = (Df4pw6 & Kf4pw6);
assign Kf4pw6 = (~(Jo4ju6 & vis_r14_o[30]));
assign Df4pw6 = (Rf4pw6 & Yf4pw6);
assign Yf4pw6 = (~(Ep4ju6 & vis_psp_o[28]));
assign Rf4pw6 = (~(Lp4ju6 & vis_msp_o[28]));
assign Pe4pw6 = (Fg4pw6 & Mg4pw6);
assign Mg4pw6 = (~(Gq4ju6 & vis_r12_o[30]));
assign Fg4pw6 = (~(Nq4ju6 & vis_r11_o[30]));
assign Be4pw6 = (Tg4pw6 & Ah4pw6);
assign Ah4pw6 = (Hh4pw6 & Oh4pw6);
assign Oh4pw6 = (~(Wr4ju6 & vis_r10_o[30]));
assign Hh4pw6 = (~(Ds4ju6 & vis_r9_o[30]));
assign Tg4pw6 = (Y50iu6 & Vh4pw6);
assign Vh4pw6 = (~(Rs4ju6 & vis_r8_o[30]));
assign Y50iu6 = (Ci4pw6 & Ji4pw6);
assign Ji4pw6 = (Qi4pw6 & Xi4pw6);
assign Xi4pw6 = (Ej4pw6 & Lj4pw6);
assign Lj4pw6 = (~(V6now6 & vis_r2_o[30]));
assign Ej4pw6 = (~(C7now6 & vis_r6_o[30]));
assign Qi4pw6 = (Sj4pw6 & Zj4pw6);
assign Zj4pw6 = (~(X7now6 & vis_r5_o[30]));
assign Sj4pw6 = (~(E8now6 & vis_r4_o[30]));
assign Ci4pw6 = (Gk4pw6 & Nk4pw6);
assign Nk4pw6 = (Uk4pw6 & Bl4pw6);
assign Bl4pw6 = (~(N9now6 & vis_r1_o[30]));
assign Uk4pw6 = (~(U9now6 & vis_r0_o[30]));
assign Gk4pw6 = (Il4pw6 & Pl4pw6);
assign Pl4pw6 = (~(Panow6 & vis_r3_o[30]));
assign Il4pw6 = (~(Wanow6 & vis_r7_o[30]));
assign Galiu6 = (!Fkfpw6[30]);
assign Gd4pw6 = (Wl4pw6 & Dm4pw6);
assign Dm4pw6 = (~(Eafpw6[30] & A3iiu6));
assign Wl4pw6 = (~(N5fpw6[29] & Sdaiu6));
assign HADDR[29] = (Xg6iu6 ? Jshpw6[29] : Dx0iu6);
assign Xg6iu6 = (!Ze9iu6);
assign Dx0iu6 = (~(Km4pw6 & Rm4pw6));
assign Rm4pw6 = (T2iiu6 | Pi0iu6);
assign Pi0iu6 = (Mm4ju6 ? Ym4pw6 : Sm8iu6);
assign Ym4pw6 = (Fn4pw6 & Mn4pw6);
assign Mn4pw6 = (Tn4pw6 & Ao4pw6);
assign Ao4pw6 = (Ho4pw6 & Oo4pw6);
assign Oo4pw6 = (~(Jo4ju6 & vis_r14_o[29]));
assign Ho4pw6 = (Vo4pw6 & Cp4pw6);
assign Cp4pw6 = (~(Ep4ju6 & vis_psp_o[27]));
assign Vo4pw6 = (~(Lp4ju6 & vis_msp_o[27]));
assign Tn4pw6 = (Jp4pw6 & Qp4pw6);
assign Qp4pw6 = (~(Gq4ju6 & vis_r12_o[29]));
assign Jp4pw6 = (~(Nq4ju6 & vis_r11_o[29]));
assign Fn4pw6 = (Xp4pw6 & Eq4pw6);
assign Eq4pw6 = (Lq4pw6 & Sq4pw6);
assign Sq4pw6 = (~(Wr4ju6 & vis_r10_o[29]));
assign Lq4pw6 = (~(Ds4ju6 & vis_r9_o[29]));
assign Xp4pw6 = (M60iu6 & Zq4pw6);
assign Zq4pw6 = (~(Rs4ju6 & vis_r8_o[29]));
assign M60iu6 = (Gr4pw6 & Nr4pw6);
assign Nr4pw6 = (Ur4pw6 & Bs4pw6);
assign Bs4pw6 = (Is4pw6 & Ps4pw6);
assign Ps4pw6 = (~(V6now6 & vis_r2_o[29]));
assign Is4pw6 = (~(C7now6 & vis_r6_o[29]));
assign Ur4pw6 = (Ws4pw6 & Dt4pw6);
assign Dt4pw6 = (~(X7now6 & vis_r5_o[29]));
assign Ws4pw6 = (~(E8now6 & vis_r4_o[29]));
assign Gr4pw6 = (Kt4pw6 & Rt4pw6);
assign Rt4pw6 = (Yt4pw6 & Fu4pw6);
assign Fu4pw6 = (~(N9now6 & vis_r1_o[29]));
assign Yt4pw6 = (~(U9now6 & vis_r0_o[29]));
assign Kt4pw6 = (Mu4pw6 & Tu4pw6);
assign Tu4pw6 = (~(Panow6 & vis_r3_o[29]));
assign Mu4pw6 = (~(Wanow6 & vis_r7_o[29]));
assign Sm8iu6 = (!Fkfpw6[29]);
assign Km4pw6 = (Av4pw6 & Hv4pw6);
assign Hv4pw6 = (~(Eafpw6[29] & A3iiu6));
assign Av4pw6 = (~(N5fpw6[28] & Sdaiu6));
assign HADDR[28] = (Ze9iu6 ? V0epw6 : Jshpw6[28]);
assign V0epw6 = (~(Ov4pw6 & Vv4pw6));
assign Vv4pw6 = (T2iiu6 | Wi0iu6);
assign Wi0iu6 = (Mm4ju6 ? Cw4pw6 : Seniu6);
assign Cw4pw6 = (Jw4pw6 & Qw4pw6);
assign Qw4pw6 = (Xw4pw6 & Ex4pw6);
assign Ex4pw6 = (Lx4pw6 & Sx4pw6);
assign Sx4pw6 = (~(Jo4ju6 & vis_r14_o[28]));
assign Lx4pw6 = (Zx4pw6 & Gy4pw6);
assign Gy4pw6 = (~(Ep4ju6 & vis_psp_o[26]));
assign Zx4pw6 = (~(Lp4ju6 & vis_msp_o[26]));
assign Xw4pw6 = (Ny4pw6 & Uy4pw6);
assign Uy4pw6 = (~(Gq4ju6 & vis_r12_o[28]));
assign Ny4pw6 = (~(Nq4ju6 & vis_r11_o[28]));
assign Jw4pw6 = (Bz4pw6 & Iz4pw6);
assign Iz4pw6 = (Pz4pw6 & Wz4pw6);
assign Wz4pw6 = (~(Wr4ju6 & vis_r10_o[28]));
assign Pz4pw6 = (~(Ds4ju6 & vis_r9_o[28]));
assign Bz4pw6 = (T60iu6 & D05pw6);
assign D05pw6 = (~(Rs4ju6 & vis_r8_o[28]));
assign T60iu6 = (!Ltnow6);
assign Ltnow6 = (~(K05pw6 & R05pw6));
assign R05pw6 = (Y05pw6 & F15pw6);
assign F15pw6 = (M15pw6 & T15pw6);
assign T15pw6 = (~(V6now6 & vis_r2_o[28]));
assign M15pw6 = (~(C7now6 & vis_r6_o[28]));
assign Y05pw6 = (A25pw6 & H25pw6);
assign H25pw6 = (~(X7now6 & vis_r5_o[28]));
assign A25pw6 = (~(E8now6 & vis_r4_o[28]));
assign K05pw6 = (O25pw6 & V25pw6);
assign V25pw6 = (C35pw6 & J35pw6);
assign J35pw6 = (~(N9now6 & vis_r1_o[28]));
assign C35pw6 = (~(U9now6 & vis_r0_o[28]));
assign O25pw6 = (Q35pw6 & X35pw6);
assign X35pw6 = (~(Panow6 & vis_r3_o[28]));
assign Q35pw6 = (~(Wanow6 & vis_r7_o[28]));
assign Seniu6 = (!Fkfpw6[28]);
assign Ov4pw6 = (E45pw6 & L45pw6);
assign L45pw6 = (~(N5fpw6[27] & Sdaiu6));
assign E45pw6 = (~(Eafpw6[28] & A3iiu6));
assign HADDR[27] = (Ze9iu6 ? O0epw6 : Jshpw6[27]);
assign O0epw6 = (~(S45pw6 & Z45pw6));
assign Z45pw6 = (~(B7iiu6 & Dj0iu6));
assign Dj0iu6 = (Cn5ju6 ? Fkfpw6[27] : G55pw6);
assign G55pw6 = (~(N55pw6 & U55pw6));
assign U55pw6 = (B65pw6 & I65pw6);
assign I65pw6 = (P65pw6 & W65pw6);
assign W65pw6 = (~(Jo4ju6 & vis_r14_o[27]));
assign P65pw6 = (D75pw6 & K75pw6);
assign K75pw6 = (~(Ep4ju6 & vis_psp_o[25]));
assign D75pw6 = (~(Lp4ju6 & vis_msp_o[25]));
assign B65pw6 = (R75pw6 & Y75pw6);
assign Y75pw6 = (~(Gq4ju6 & vis_r12_o[27]));
assign R75pw6 = (~(Nq4ju6 & vis_r11_o[27]));
assign N55pw6 = (F85pw6 & M85pw6);
assign M85pw6 = (T85pw6 & A95pw6);
assign A95pw6 = (~(Wr4ju6 & vis_r10_o[27]));
assign T85pw6 = (~(Ds4ju6 & vis_r9_o[27]));
assign F85pw6 = (A70iu6 & H95pw6);
assign H95pw6 = (~(Rs4ju6 & vis_r8_o[27]));
assign A70iu6 = (O95pw6 & V95pw6);
assign V95pw6 = (Ca5pw6 & Ja5pw6);
assign Ja5pw6 = (Qa5pw6 & Xa5pw6);
assign Xa5pw6 = (~(V6now6 & vis_r2_o[27]));
assign Qa5pw6 = (~(C7now6 & vis_r6_o[27]));
assign Ca5pw6 = (Eb5pw6 & Lb5pw6);
assign Lb5pw6 = (~(X7now6 & vis_r5_o[27]));
assign Eb5pw6 = (~(E8now6 & vis_r4_o[27]));
assign O95pw6 = (Sb5pw6 & Zb5pw6);
assign Zb5pw6 = (Gc5pw6 & Nc5pw6);
assign Nc5pw6 = (~(N9now6 & vis_r1_o[27]));
assign Gc5pw6 = (~(U9now6 & vis_r0_o[27]));
assign Sb5pw6 = (Uc5pw6 & Bd5pw6);
assign Bd5pw6 = (~(Panow6 & vis_r3_o[27]));
assign Uc5pw6 = (~(Wanow6 & vis_r7_o[27]));
assign S45pw6 = (Id5pw6 & Pd5pw6);
assign Pd5pw6 = (~(N5fpw6[26] & Sdaiu6));
assign Id5pw6 = (~(Eafpw6[27] & A3iiu6));
assign HADDR[26] = (Ze9iu6 ? H0epw6 : Jshpw6[26]);
assign H0epw6 = (~(Wd5pw6 & De5pw6));
assign De5pw6 = (~(B7iiu6 & Kj0iu6));
assign Kj0iu6 = (Cn5ju6 ? Fkfpw6[26] : Ke5pw6);
assign Ke5pw6 = (~(Re5pw6 & Ye5pw6));
assign Ye5pw6 = (Ff5pw6 & Mf5pw6);
assign Mf5pw6 = (Tf5pw6 & Ag5pw6);
assign Ag5pw6 = (~(Jo4ju6 & vis_r14_o[26]));
assign Tf5pw6 = (Hg5pw6 & Og5pw6);
assign Og5pw6 = (~(Ep4ju6 & vis_psp_o[24]));
assign Hg5pw6 = (~(Lp4ju6 & vis_msp_o[24]));
assign Ff5pw6 = (Vg5pw6 & Ch5pw6);
assign Ch5pw6 = (~(Gq4ju6 & vis_r12_o[26]));
assign Vg5pw6 = (~(Nq4ju6 & vis_r11_o[26]));
assign Re5pw6 = (Jh5pw6 & Qh5pw6);
assign Qh5pw6 = (Xh5pw6 & Ei5pw6);
assign Ei5pw6 = (~(Wr4ju6 & vis_r10_o[26]));
assign Xh5pw6 = (~(Ds4ju6 & vis_r9_o[26]));
assign Jh5pw6 = (H70iu6 & Li5pw6);
assign Li5pw6 = (~(Rs4ju6 & vis_r8_o[26]));
assign H70iu6 = (Si5pw6 & Zi5pw6);
assign Zi5pw6 = (Gj5pw6 & Nj5pw6);
assign Nj5pw6 = (Uj5pw6 & Bk5pw6);
assign Bk5pw6 = (~(V6now6 & vis_r2_o[26]));
assign Uj5pw6 = (~(C7now6 & vis_r6_o[26]));
assign Gj5pw6 = (Ik5pw6 & Pk5pw6);
assign Pk5pw6 = (~(X7now6 & vis_r5_o[26]));
assign Ik5pw6 = (~(E8now6 & vis_r4_o[26]));
assign Si5pw6 = (Wk5pw6 & Dl5pw6);
assign Dl5pw6 = (Kl5pw6 & Rl5pw6);
assign Rl5pw6 = (~(N9now6 & vis_r1_o[26]));
assign Kl5pw6 = (~(U9now6 & vis_r0_o[26]));
assign Wk5pw6 = (Yl5pw6 & Fm5pw6);
assign Fm5pw6 = (~(Panow6 & vis_r3_o[26]));
assign Yl5pw6 = (~(Wanow6 & vis_r7_o[26]));
assign Wd5pw6 = (Mm5pw6 & Tm5pw6);
assign Tm5pw6 = (~(N5fpw6[25] & Sdaiu6));
assign Mm5pw6 = (~(Eafpw6[26] & A3iiu6));
assign HADDR[25] = (Ze9iu6 ? A0epw6 : Jshpw6[25]);
assign A0epw6 = (~(An5pw6 & Hn5pw6));
assign Hn5pw6 = (~(B7iiu6 & Rj0iu6));
assign Rj0iu6 = (Cn5ju6 ? Fkfpw6[25] : On5pw6);
assign On5pw6 = (~(Vn5pw6 & Co5pw6));
assign Co5pw6 = (Jo5pw6 & Qo5pw6);
assign Qo5pw6 = (Xo5pw6 & Ep5pw6);
assign Ep5pw6 = (~(Jo4ju6 & vis_r14_o[25]));
assign Xo5pw6 = (Lp5pw6 & Sp5pw6);
assign Sp5pw6 = (~(Ep4ju6 & vis_psp_o[23]));
assign Lp5pw6 = (~(Lp4ju6 & vis_msp_o[23]));
assign Jo5pw6 = (Zp5pw6 & Gq5pw6);
assign Gq5pw6 = (~(Gq4ju6 & vis_r12_o[25]));
assign Zp5pw6 = (~(Nq4ju6 & vis_r11_o[25]));
assign Vn5pw6 = (Nq5pw6 & Uq5pw6);
assign Uq5pw6 = (Br5pw6 & Ir5pw6);
assign Ir5pw6 = (~(Wr4ju6 & vis_r10_o[25]));
assign Br5pw6 = (~(Ds4ju6 & vis_r9_o[25]));
assign Nq5pw6 = (O70iu6 & Pr5pw6);
assign Pr5pw6 = (~(Rs4ju6 & vis_r8_o[25]));
assign O70iu6 = (Wr5pw6 & Ds5pw6);
assign Ds5pw6 = (Ks5pw6 & Rs5pw6);
assign Rs5pw6 = (Ys5pw6 & Ft5pw6);
assign Ft5pw6 = (~(V6now6 & vis_r2_o[25]));
assign Ys5pw6 = (~(C7now6 & vis_r6_o[25]));
assign Ks5pw6 = (Mt5pw6 & Tt5pw6);
assign Tt5pw6 = (~(X7now6 & vis_r5_o[25]));
assign Mt5pw6 = (~(E8now6 & vis_r4_o[25]));
assign Wr5pw6 = (Au5pw6 & Hu5pw6);
assign Hu5pw6 = (Ou5pw6 & Vu5pw6);
assign Vu5pw6 = (~(N9now6 & vis_r1_o[25]));
assign Ou5pw6 = (~(U9now6 & vis_r0_o[25]));
assign Au5pw6 = (Cv5pw6 & Jv5pw6);
assign Jv5pw6 = (~(Panow6 & vis_r3_o[25]));
assign Cv5pw6 = (~(Wanow6 & vis_r7_o[25]));
assign An5pw6 = (Qv5pw6 & Xv5pw6);
assign Xv5pw6 = (~(N5fpw6[24] & Sdaiu6));
assign Qv5pw6 = (~(Eafpw6[25] & A3iiu6));
assign HADDR[24] = (Ze9iu6 ? Tzdpw6 : Jshpw6[24]);
assign Tzdpw6 = (~(Ew5pw6 & Lw5pw6));
assign Lw5pw6 = (T2iiu6 | Yj0iu6);
assign Yj0iu6 = (Mm4ju6 ? Sw5pw6 : Kykiu6);
assign Sw5pw6 = (Zw5pw6 & Gx5pw6);
assign Gx5pw6 = (Nx5pw6 & Ux5pw6);
assign Ux5pw6 = (By5pw6 & Iy5pw6);
assign Iy5pw6 = (~(Jo4ju6 & vis_r14_o[24]));
assign By5pw6 = (Py5pw6 & Wy5pw6);
assign Wy5pw6 = (~(Ep4ju6 & vis_psp_o[22]));
assign Py5pw6 = (~(Lp4ju6 & vis_msp_o[22]));
assign Nx5pw6 = (Dz5pw6 & Kz5pw6);
assign Kz5pw6 = (~(Gq4ju6 & vis_r12_o[24]));
assign Dz5pw6 = (~(Nq4ju6 & vis_r11_o[24]));
assign Zw5pw6 = (Rz5pw6 & Yz5pw6);
assign Yz5pw6 = (F06pw6 & M06pw6);
assign M06pw6 = (~(Wr4ju6 & vis_r10_o[24]));
assign F06pw6 = (~(Ds4ju6 & vis_r9_o[24]));
assign Rz5pw6 = (V70iu6 & T06pw6);
assign T06pw6 = (~(Rs4ju6 & vis_r8_o[24]));
assign V70iu6 = (A16pw6 & H16pw6);
assign H16pw6 = (O16pw6 & V16pw6);
assign V16pw6 = (C26pw6 & J26pw6);
assign J26pw6 = (~(V6now6 & vis_r2_o[24]));
assign C26pw6 = (~(C7now6 & vis_r6_o[24]));
assign O16pw6 = (Q26pw6 & X26pw6);
assign X26pw6 = (~(X7now6 & vis_r5_o[24]));
assign Q26pw6 = (~(E8now6 & vis_r4_o[24]));
assign A16pw6 = (E36pw6 & L36pw6);
assign L36pw6 = (S36pw6 & Z36pw6);
assign Z36pw6 = (~(N9now6 & vis_r1_o[24]));
assign S36pw6 = (~(U9now6 & vis_r0_o[24]));
assign E36pw6 = (G46pw6 & N46pw6);
assign N46pw6 = (~(Panow6 & vis_r3_o[24]));
assign G46pw6 = (~(Wanow6 & vis_r7_o[24]));
assign Kykiu6 = (!Fkfpw6[24]);
assign Ew5pw6 = (U46pw6 & B56pw6);
assign B56pw6 = (~(N5fpw6[23] & Sdaiu6));
assign U46pw6 = (~(Eafpw6[24] & A3iiu6));
assign HADDR[23] = (Ze9iu6 ? Mzdpw6 : Jshpw6[23]);
assign Mzdpw6 = (~(I56pw6 & P56pw6));
assign P56pw6 = (T2iiu6 | Fk0iu6);
assign Fk0iu6 = (Mm4ju6 ? W56pw6 : Ax9iu6);
assign W56pw6 = (D66pw6 & K66pw6);
assign K66pw6 = (R66pw6 & Y66pw6);
assign Y66pw6 = (F76pw6 & M76pw6);
assign M76pw6 = (~(Jo4ju6 & vis_r14_o[23]));
assign F76pw6 = (T76pw6 & A86pw6);
assign A86pw6 = (~(Ep4ju6 & vis_psp_o[21]));
assign T76pw6 = (~(Lp4ju6 & vis_msp_o[21]));
assign R66pw6 = (H86pw6 & O86pw6);
assign O86pw6 = (~(Gq4ju6 & vis_r12_o[23]));
assign H86pw6 = (~(Nq4ju6 & vis_r11_o[23]));
assign D66pw6 = (V86pw6 & C96pw6);
assign C96pw6 = (J96pw6 & Q96pw6);
assign Q96pw6 = (~(Wr4ju6 & vis_r10_o[23]));
assign J96pw6 = (~(Ds4ju6 & vis_r9_o[23]));
assign V86pw6 = (C80iu6 & X96pw6);
assign X96pw6 = (~(Rs4ju6 & vis_r8_o[23]));
assign C80iu6 = (Ea6pw6 & La6pw6);
assign La6pw6 = (Sa6pw6 & Za6pw6);
assign Za6pw6 = (Gb6pw6 & Nb6pw6);
assign Nb6pw6 = (~(V6now6 & vis_r2_o[23]));
assign Gb6pw6 = (~(C7now6 & vis_r6_o[23]));
assign Sa6pw6 = (Ub6pw6 & Bc6pw6);
assign Bc6pw6 = (~(X7now6 & vis_r5_o[23]));
assign Ub6pw6 = (~(E8now6 & vis_r4_o[23]));
assign Ea6pw6 = (Ic6pw6 & Pc6pw6);
assign Pc6pw6 = (Wc6pw6 & Dd6pw6);
assign Dd6pw6 = (~(N9now6 & vis_r1_o[23]));
assign Wc6pw6 = (~(U9now6 & vis_r0_o[23]));
assign Ic6pw6 = (Kd6pw6 & Rd6pw6);
assign Rd6pw6 = (~(Panow6 & vis_r3_o[23]));
assign Kd6pw6 = (~(Wanow6 & vis_r7_o[23]));
assign Ax9iu6 = (!Fkfpw6[23]);
assign I56pw6 = (Yd6pw6 & Fe6pw6);
assign Fe6pw6 = (~(N5fpw6[22] & Sdaiu6));
assign Yd6pw6 = (~(Eafpw6[23] & A3iiu6));
assign HADDR[22] = (Ze9iu6 ? Fzdpw6 : Jshpw6[22]);
assign Fzdpw6 = (~(Me6pw6 & Te6pw6));
assign Te6pw6 = (T2iiu6 | Mk0iu6);
assign Mk0iu6 = (Mm4ju6 ? Af6pw6 : Suliu6);
assign Af6pw6 = (Hf6pw6 & Of6pw6);
assign Of6pw6 = (Vf6pw6 & Cg6pw6);
assign Cg6pw6 = (Jg6pw6 & Qg6pw6);
assign Qg6pw6 = (~(Jo4ju6 & vis_r14_o[22]));
assign Jg6pw6 = (Xg6pw6 & Eh6pw6);
assign Eh6pw6 = (~(Ep4ju6 & vis_psp_o[20]));
assign Xg6pw6 = (~(Lp4ju6 & vis_msp_o[20]));
assign Vf6pw6 = (Lh6pw6 & Sh6pw6);
assign Sh6pw6 = (~(Gq4ju6 & vis_r12_o[22]));
assign Lh6pw6 = (~(Nq4ju6 & vis_r11_o[22]));
assign Hf6pw6 = (Zh6pw6 & Gi6pw6);
assign Gi6pw6 = (Ni6pw6 & Ui6pw6);
assign Ui6pw6 = (~(Wr4ju6 & vis_r10_o[22]));
assign Ni6pw6 = (~(Ds4ju6 & vis_r9_o[22]));
assign Zh6pw6 = (J80iu6 & Bj6pw6);
assign Bj6pw6 = (~(Rs4ju6 & vis_r8_o[22]));
assign J80iu6 = (Ij6pw6 & Pj6pw6);
assign Pj6pw6 = (Wj6pw6 & Dk6pw6);
assign Dk6pw6 = (Kk6pw6 & Rk6pw6);
assign Rk6pw6 = (~(V6now6 & vis_r2_o[22]));
assign Kk6pw6 = (~(C7now6 & vis_r6_o[22]));
assign Wj6pw6 = (Yk6pw6 & Fl6pw6);
assign Fl6pw6 = (~(X7now6 & vis_r5_o[22]));
assign Yk6pw6 = (~(E8now6 & vis_r4_o[22]));
assign Ij6pw6 = (Ml6pw6 & Tl6pw6);
assign Tl6pw6 = (Am6pw6 & Hm6pw6);
assign Hm6pw6 = (~(N9now6 & vis_r1_o[22]));
assign Am6pw6 = (~(U9now6 & vis_r0_o[22]));
assign Ml6pw6 = (Om6pw6 & Vm6pw6);
assign Vm6pw6 = (~(Panow6 & vis_r3_o[22]));
assign Om6pw6 = (~(Wanow6 & vis_r7_o[22]));
assign Suliu6 = (!Fkfpw6[22]);
assign Me6pw6 = (Cn6pw6 & Jn6pw6);
assign Jn6pw6 = (~(N5fpw6[21] & Sdaiu6));
assign Cn6pw6 = (~(Eafpw6[22] & A3iiu6));
assign HADDR[21] = (Ze9iu6 ? Yydpw6 : Jshpw6[21]);
assign Yydpw6 = (~(Qn6pw6 & Xn6pw6));
assign Xn6pw6 = (T2iiu6 | Tk0iu6);
assign Tk0iu6 = (Mm4ju6 ? Eo6pw6 : Rxliu6);
assign Eo6pw6 = (Lo6pw6 & So6pw6);
assign So6pw6 = (Zo6pw6 & Gp6pw6);
assign Gp6pw6 = (Np6pw6 & Up6pw6);
assign Up6pw6 = (~(Jo4ju6 & vis_r14_o[21]));
assign Np6pw6 = (Bq6pw6 & Iq6pw6);
assign Iq6pw6 = (~(Ep4ju6 & vis_psp_o[19]));
assign Bq6pw6 = (~(Lp4ju6 & vis_msp_o[19]));
assign Zo6pw6 = (Pq6pw6 & Wq6pw6);
assign Wq6pw6 = (~(Gq4ju6 & vis_r12_o[21]));
assign Pq6pw6 = (~(Nq4ju6 & vis_r11_o[21]));
assign Lo6pw6 = (Dr6pw6 & Kr6pw6);
assign Kr6pw6 = (Rr6pw6 & Yr6pw6);
assign Yr6pw6 = (~(Wr4ju6 & vis_r10_o[21]));
assign Rr6pw6 = (~(Ds4ju6 & vis_r9_o[21]));
assign Dr6pw6 = (Q80iu6 & Fs6pw6);
assign Fs6pw6 = (~(Rs4ju6 & vis_r8_o[21]));
assign Q80iu6 = (Ms6pw6 & Ts6pw6);
assign Ts6pw6 = (At6pw6 & Ht6pw6);
assign Ht6pw6 = (Ot6pw6 & Vt6pw6);
assign Vt6pw6 = (~(V6now6 & vis_r2_o[21]));
assign Ot6pw6 = (~(C7now6 & vis_r6_o[21]));
assign At6pw6 = (Cu6pw6 & Ju6pw6);
assign Ju6pw6 = (~(X7now6 & vis_r5_o[21]));
assign Cu6pw6 = (~(E8now6 & vis_r4_o[21]));
assign Ms6pw6 = (Qu6pw6 & Xu6pw6);
assign Xu6pw6 = (Ev6pw6 & Lv6pw6);
assign Lv6pw6 = (~(N9now6 & vis_r1_o[21]));
assign Ev6pw6 = (~(U9now6 & vis_r0_o[21]));
assign Qu6pw6 = (Sv6pw6 & Zv6pw6);
assign Zv6pw6 = (~(Panow6 & vis_r3_o[21]));
assign Sv6pw6 = (~(Wanow6 & vis_r7_o[21]));
assign Rxliu6 = (!Fkfpw6[21]);
assign Qn6pw6 = (Gw6pw6 & Nw6pw6);
assign Nw6pw6 = (~(N5fpw6[20] & Sdaiu6));
assign Gw6pw6 = (~(Eafpw6[21] & A3iiu6));
assign HADDR[20] = (Ze9iu6 ? Rydpw6 : Jshpw6[20]);
assign Rydpw6 = (~(Uw6pw6 & Bx6pw6));
assign Bx6pw6 = (T2iiu6 | Al0iu6);
assign Al0iu6 = (Mm4ju6 ? Ix6pw6 : X0miu6);
assign Ix6pw6 = (Px6pw6 & Wx6pw6);
assign Wx6pw6 = (Dy6pw6 & Ky6pw6);
assign Ky6pw6 = (Ry6pw6 & Yy6pw6);
assign Yy6pw6 = (~(Jo4ju6 & vis_r14_o[20]));
assign Ry6pw6 = (Fz6pw6 & Mz6pw6);
assign Mz6pw6 = (~(Ep4ju6 & vis_psp_o[18]));
assign Fz6pw6 = (~(Lp4ju6 & vis_msp_o[18]));
assign Dy6pw6 = (Tz6pw6 & A07pw6);
assign A07pw6 = (~(Gq4ju6 & vis_r12_o[20]));
assign Tz6pw6 = (~(Nq4ju6 & vis_r11_o[20]));
assign Px6pw6 = (H07pw6 & O07pw6);
assign O07pw6 = (V07pw6 & C17pw6);
assign C17pw6 = (~(Wr4ju6 & vis_r10_o[20]));
assign V07pw6 = (~(Ds4ju6 & vis_r9_o[20]));
assign H07pw6 = (X80iu6 & J17pw6);
assign J17pw6 = (~(Rs4ju6 & vis_r8_o[20]));
assign X80iu6 = (Q17pw6 & X17pw6);
assign X17pw6 = (E27pw6 & L27pw6);
assign L27pw6 = (S27pw6 & Z27pw6);
assign Z27pw6 = (~(V6now6 & vis_r2_o[20]));
assign S27pw6 = (~(C7now6 & vis_r6_o[20]));
assign E27pw6 = (G37pw6 & N37pw6);
assign N37pw6 = (~(X7now6 & vis_r5_o[20]));
assign G37pw6 = (~(E8now6 & vis_r4_o[20]));
assign Q17pw6 = (U37pw6 & B47pw6);
assign B47pw6 = (I47pw6 & P47pw6);
assign P47pw6 = (~(N9now6 & vis_r1_o[20]));
assign I47pw6 = (~(U9now6 & vis_r0_o[20]));
assign U37pw6 = (W47pw6 & D57pw6);
assign D57pw6 = (~(Panow6 & vis_r3_o[20]));
assign W47pw6 = (~(Wanow6 & vis_r7_o[20]));
assign X0miu6 = (!Fkfpw6[20]);
assign Uw6pw6 = (K57pw6 & R57pw6);
assign R57pw6 = (~(N5fpw6[19] & Sdaiu6));
assign K57pw6 = (~(Eafpw6[20] & A3iiu6));
assign HADDR[1] = (~(Y57pw6 & F67pw6));
assign F67pw6 = (~(M67pw6 & Ne3pw6));
assign M67pw6 = (Tnhpw6[1] & T67pw6);
assign T67pw6 = (!Aphpw6[2]);
assign Y57pw6 = (~(Hz0iu6 & Ze9iu6));
assign Hz0iu6 = (A77pw6 & Ed3pw6);
assign A77pw6 = (Iiliu6 & Ob3pw6);
assign Iiliu6 = (~(H77pw6 & O77pw6));
assign O77pw6 = (T2iiu6 | Hl0iu6);
assign Hl0iu6 = (Mm4ju6 ? V77pw6 : Rjliu6);
assign V77pw6 = (C87pw6 & J87pw6);
assign J87pw6 = (Q87pw6 & X87pw6);
assign X87pw6 = (E97pw6 & L97pw6);
assign L97pw6 = (~(Jo4ju6 & vis_r14_o[1]));
assign E97pw6 = (~(Gq4ju6 & vis_r12_o[1]));
assign Q87pw6 = (S97pw6 & Z97pw6);
assign Z97pw6 = (~(Nq4ju6 & vis_r11_o[1]));
assign S97pw6 = (~(Wr4ju6 & vis_r10_o[1]));
assign C87pw6 = (Ga7pw6 & E90iu6);
assign E90iu6 = (Na7pw6 & Ua7pw6);
assign Ua7pw6 = (Bb7pw6 & Ib7pw6);
assign Ib7pw6 = (Pb7pw6 & Wb7pw6);
assign Wb7pw6 = (~(V6now6 & vis_r2_o[1]));
assign Pb7pw6 = (~(C7now6 & vis_r6_o[1]));
assign Bb7pw6 = (Dc7pw6 & Kc7pw6);
assign Kc7pw6 = (~(X7now6 & vis_r5_o[1]));
assign Dc7pw6 = (~(E8now6 & vis_r4_o[1]));
assign Na7pw6 = (Rc7pw6 & Yc7pw6);
assign Yc7pw6 = (Fd7pw6 & Md7pw6);
assign Md7pw6 = (~(N9now6 & vis_r1_o[1]));
assign Fd7pw6 = (~(U9now6 & vis_r0_o[1]));
assign Rc7pw6 = (Td7pw6 & Ae7pw6);
assign Ae7pw6 = (~(Panow6 & vis_r3_o[1]));
assign Td7pw6 = (~(Wanow6 & vis_r7_o[1]));
assign Ga7pw6 = (He7pw6 & Oe7pw6);
assign Oe7pw6 = (~(Ds4ju6 & vis_r9_o[1]));
assign He7pw6 = (~(Rs4ju6 & vis_r8_o[1]));
assign Rjliu6 = (!Fkfpw6[1]);
assign H77pw6 = (Ve7pw6 & Cf7pw6);
assign Cf7pw6 = (~(Jf7pw6 & Sdaiu6));
assign Jf7pw6 = (~(Qf7pw6 | Vtzhu6));
assign Vtzhu6 = (Pkciu6 & vis_pc_o[0]);
assign Qf7pw6 = (~(Pkciu6 | vis_pc_o[0]));
assign Ve7pw6 = (~(Eafpw6[1] & A3iiu6));
assign HADDR[19] = (Ze9iu6 ? Kydpw6 : Jshpw6[19]);
assign Kydpw6 = (~(Xf7pw6 & Eg7pw6));
assign Eg7pw6 = (T2iiu6 | Ol0iu6);
assign Ol0iu6 = (Mm4ju6 ? Lg7pw6 : W3miu6);
assign Lg7pw6 = (Sg7pw6 & Zg7pw6);
assign Zg7pw6 = (Gh7pw6 & Nh7pw6);
assign Nh7pw6 = (Uh7pw6 & Bi7pw6);
assign Bi7pw6 = (~(Jo4ju6 & vis_r14_o[19]));
assign Uh7pw6 = (Ii7pw6 & Pi7pw6);
assign Pi7pw6 = (~(Ep4ju6 & vis_psp_o[17]));
assign Ii7pw6 = (~(Lp4ju6 & vis_msp_o[17]));
assign Gh7pw6 = (Wi7pw6 & Dj7pw6);
assign Dj7pw6 = (~(Gq4ju6 & vis_r12_o[19]));
assign Wi7pw6 = (~(Nq4ju6 & vis_r11_o[19]));
assign Sg7pw6 = (Kj7pw6 & Rj7pw6);
assign Rj7pw6 = (Yj7pw6 & Fk7pw6);
assign Fk7pw6 = (~(Wr4ju6 & vis_r10_o[19]));
assign Yj7pw6 = (~(Ds4ju6 & vis_r9_o[19]));
assign Kj7pw6 = (L90iu6 & Mk7pw6);
assign Mk7pw6 = (~(Rs4ju6 & vis_r8_o[19]));
assign L90iu6 = (Tk7pw6 & Al7pw6);
assign Al7pw6 = (Hl7pw6 & Ol7pw6);
assign Ol7pw6 = (Vl7pw6 & Cm7pw6);
assign Cm7pw6 = (~(V6now6 & vis_r2_o[19]));
assign Vl7pw6 = (~(C7now6 & vis_r6_o[19]));
assign Hl7pw6 = (Jm7pw6 & Qm7pw6);
assign Qm7pw6 = (~(X7now6 & vis_r5_o[19]));
assign Jm7pw6 = (~(E8now6 & vis_r4_o[19]));
assign Tk7pw6 = (Xm7pw6 & En7pw6);
assign En7pw6 = (Ln7pw6 & Sn7pw6);
assign Sn7pw6 = (~(N9now6 & vis_r1_o[19]));
assign Ln7pw6 = (~(U9now6 & vis_r0_o[19]));
assign Xm7pw6 = (Zn7pw6 & Go7pw6);
assign Go7pw6 = (~(Panow6 & vis_r3_o[19]));
assign Zn7pw6 = (~(Wanow6 & vis_r7_o[19]));
assign W3miu6 = (!Fkfpw6[19]);
assign Xf7pw6 = (No7pw6 & Uo7pw6);
assign Uo7pw6 = (~(N5fpw6[18] & Sdaiu6));
assign No7pw6 = (~(Eafpw6[19] & A3iiu6));
assign HADDR[18] = (Ze9iu6 ? Dydpw6 : Jshpw6[18]);
assign Dydpw6 = (~(Bp7pw6 & Ip7pw6));
assign Ip7pw6 = (T2iiu6 | Vl0iu6);
assign Vl0iu6 = (Mm4ju6 ? Pp7pw6 : V6miu6);
assign Pp7pw6 = (Wp7pw6 & Dq7pw6);
assign Dq7pw6 = (Kq7pw6 & Rq7pw6);
assign Rq7pw6 = (Yq7pw6 & Fr7pw6);
assign Fr7pw6 = (~(Jo4ju6 & vis_r14_o[18]));
assign Yq7pw6 = (Mr7pw6 & Tr7pw6);
assign Tr7pw6 = (~(Ep4ju6 & vis_psp_o[16]));
assign Mr7pw6 = (~(Lp4ju6 & vis_msp_o[16]));
assign Kq7pw6 = (As7pw6 & Hs7pw6);
assign Hs7pw6 = (~(Gq4ju6 & vis_r12_o[18]));
assign As7pw6 = (~(Nq4ju6 & vis_r11_o[18]));
assign Wp7pw6 = (Os7pw6 & Vs7pw6);
assign Vs7pw6 = (Ct7pw6 & Jt7pw6);
assign Jt7pw6 = (~(Wr4ju6 & vis_r10_o[18]));
assign Ct7pw6 = (~(Ds4ju6 & vis_r9_o[18]));
assign Os7pw6 = (S90iu6 & Qt7pw6);
assign Qt7pw6 = (~(Rs4ju6 & vis_r8_o[18]));
assign S90iu6 = (Xt7pw6 & Eu7pw6);
assign Eu7pw6 = (Lu7pw6 & Su7pw6);
assign Su7pw6 = (Zu7pw6 & Gv7pw6);
assign Gv7pw6 = (~(V6now6 & vis_r2_o[18]));
assign Zu7pw6 = (~(C7now6 & vis_r6_o[18]));
assign Lu7pw6 = (Nv7pw6 & Uv7pw6);
assign Uv7pw6 = (~(X7now6 & vis_r5_o[18]));
assign Nv7pw6 = (~(E8now6 & vis_r4_o[18]));
assign Xt7pw6 = (Bw7pw6 & Iw7pw6);
assign Iw7pw6 = (Pw7pw6 & Ww7pw6);
assign Ww7pw6 = (~(N9now6 & vis_r1_o[18]));
assign Pw7pw6 = (~(U9now6 & vis_r0_o[18]));
assign Bw7pw6 = (Dx7pw6 & Kx7pw6);
assign Kx7pw6 = (~(Panow6 & vis_r3_o[18]));
assign Dx7pw6 = (~(Wanow6 & vis_r7_o[18]));
assign V6miu6 = (!Fkfpw6[18]);
assign Bp7pw6 = (Rx7pw6 & Yx7pw6);
assign Yx7pw6 = (~(N5fpw6[17] & Sdaiu6));
assign Rx7pw6 = (~(Eafpw6[18] & A3iiu6));
assign HADDR[17] = (Ze9iu6 ? Wxdpw6 : Jshpw6[17]);
assign Wxdpw6 = (~(Fy7pw6 & My7pw6));
assign My7pw6 = (T2iiu6 | Cm0iu6);
assign Cm0iu6 = (Mm4ju6 ? Ty7pw6 : U9miu6);
assign Ty7pw6 = (Az7pw6 & Hz7pw6);
assign Hz7pw6 = (Oz7pw6 & Vz7pw6);
assign Vz7pw6 = (C08pw6 & J08pw6);
assign J08pw6 = (~(Jo4ju6 & vis_r14_o[17]));
assign C08pw6 = (Q08pw6 & X08pw6);
assign X08pw6 = (~(Ep4ju6 & vis_psp_o[15]));
assign Q08pw6 = (~(Lp4ju6 & vis_msp_o[15]));
assign Oz7pw6 = (E18pw6 & L18pw6);
assign L18pw6 = (~(Gq4ju6 & vis_r12_o[17]));
assign E18pw6 = (~(Nq4ju6 & vis_r11_o[17]));
assign Az7pw6 = (S18pw6 & Z18pw6);
assign Z18pw6 = (G28pw6 & N28pw6);
assign N28pw6 = (~(Wr4ju6 & vis_r10_o[17]));
assign G28pw6 = (~(Ds4ju6 & vis_r9_o[17]));
assign S18pw6 = (Z90iu6 & U28pw6);
assign U28pw6 = (~(Rs4ju6 & vis_r8_o[17]));
assign Z90iu6 = (B38pw6 & I38pw6);
assign I38pw6 = (P38pw6 & W38pw6);
assign W38pw6 = (D48pw6 & K48pw6);
assign K48pw6 = (~(V6now6 & vis_r2_o[17]));
assign D48pw6 = (~(C7now6 & vis_r6_o[17]));
assign P38pw6 = (R48pw6 & Y48pw6);
assign Y48pw6 = (~(X7now6 & vis_r5_o[17]));
assign R48pw6 = (~(E8now6 & vis_r4_o[17]));
assign B38pw6 = (F58pw6 & M58pw6);
assign M58pw6 = (T58pw6 & A68pw6);
assign A68pw6 = (~(N9now6 & vis_r1_o[17]));
assign T58pw6 = (~(U9now6 & vis_r0_o[17]));
assign F58pw6 = (H68pw6 & O68pw6);
assign O68pw6 = (~(Panow6 & vis_r3_o[17]));
assign H68pw6 = (~(Wanow6 & vis_r7_o[17]));
assign U9miu6 = (!Fkfpw6[17]);
assign Fy7pw6 = (V68pw6 & C78pw6);
assign C78pw6 = (~(N5fpw6[16] & Sdaiu6));
assign V68pw6 = (~(Eafpw6[17] & A3iiu6));
assign HADDR[16] = (Ze9iu6 ? Pxdpw6 : Jshpw6[16]);
assign Pxdpw6 = (~(J78pw6 & Q78pw6));
assign Q78pw6 = (T2iiu6 | Jm0iu6);
assign Jm0iu6 = (Mm4ju6 ? X78pw6 : Tcmiu6);
assign X78pw6 = (E88pw6 & L88pw6);
assign L88pw6 = (S88pw6 & Z88pw6);
assign Z88pw6 = (G98pw6 & N98pw6);
assign N98pw6 = (~(Jo4ju6 & vis_r14_o[16]));
assign G98pw6 = (U98pw6 & Ba8pw6);
assign Ba8pw6 = (~(Ep4ju6 & vis_psp_o[14]));
assign U98pw6 = (~(Lp4ju6 & vis_msp_o[14]));
assign S88pw6 = (Ia8pw6 & Pa8pw6);
assign Pa8pw6 = (~(Gq4ju6 & vis_r12_o[16]));
assign Ia8pw6 = (~(Nq4ju6 & vis_r11_o[16]));
assign E88pw6 = (Wa8pw6 & Db8pw6);
assign Db8pw6 = (Kb8pw6 & Rb8pw6);
assign Rb8pw6 = (~(Wr4ju6 & vis_r10_o[16]));
assign Kb8pw6 = (~(Ds4ju6 & vis_r9_o[16]));
assign Wa8pw6 = (Ga0iu6 & Yb8pw6);
assign Yb8pw6 = (~(Rs4ju6 & vis_r8_o[16]));
assign Ga0iu6 = (Fc8pw6 & Mc8pw6);
assign Mc8pw6 = (Tc8pw6 & Ad8pw6);
assign Ad8pw6 = (Hd8pw6 & Od8pw6);
assign Od8pw6 = (~(V6now6 & vis_r2_o[16]));
assign Hd8pw6 = (~(C7now6 & vis_r6_o[16]));
assign Tc8pw6 = (Vd8pw6 & Ce8pw6);
assign Ce8pw6 = (~(X7now6 & vis_r5_o[16]));
assign Vd8pw6 = (~(E8now6 & vis_r4_o[16]));
assign Fc8pw6 = (Je8pw6 & Qe8pw6);
assign Qe8pw6 = (Xe8pw6 & Ef8pw6);
assign Ef8pw6 = (~(N9now6 & vis_r1_o[16]));
assign Xe8pw6 = (~(U9now6 & vis_r0_o[16]));
assign Je8pw6 = (Lf8pw6 & Sf8pw6);
assign Sf8pw6 = (~(Panow6 & vis_r3_o[16]));
assign Lf8pw6 = (~(Wanow6 & vis_r7_o[16]));
assign Tcmiu6 = (!Fkfpw6[16]);
assign J78pw6 = (Zf8pw6 & Gg8pw6);
assign Gg8pw6 = (~(N5fpw6[15] & Sdaiu6));
assign Zf8pw6 = (~(Eafpw6[16] & A3iiu6));
assign HADDR[15] = (Ze9iu6 ? Tugpw6[13] : Jshpw6[15]);
assign Tugpw6[13] = (~(Ng8pw6 & Ug8pw6));
assign Ug8pw6 = (~(N5fpw6[14] & Sdaiu6));
assign Ng8pw6 = (Bh8pw6 & Ih8pw6);
assign Ih8pw6 = (T2iiu6 | Qm0iu6);
assign Qm0iu6 = (Mm4ju6 ? Ph8pw6 : Sfmiu6);
assign Ph8pw6 = (Wh8pw6 & Di8pw6);
assign Di8pw6 = (Ki8pw6 & Ri8pw6);
assign Ri8pw6 = (Yi8pw6 & Fj8pw6);
assign Fj8pw6 = (~(Jo4ju6 & vis_r14_o[15]));
assign Yi8pw6 = (Mj8pw6 & Tj8pw6);
assign Tj8pw6 = (~(Ep4ju6 & vis_psp_o[13]));
assign Mj8pw6 = (~(Lp4ju6 & vis_msp_o[13]));
assign Ki8pw6 = (Ak8pw6 & Hk8pw6);
assign Hk8pw6 = (~(Gq4ju6 & vis_r12_o[15]));
assign Ak8pw6 = (~(Nq4ju6 & vis_r11_o[15]));
assign Wh8pw6 = (Ok8pw6 & Vk8pw6);
assign Vk8pw6 = (Cl8pw6 & Jl8pw6);
assign Jl8pw6 = (~(Wr4ju6 & vis_r10_o[15]));
assign Cl8pw6 = (~(Ds4ju6 & vis_r9_o[15]));
assign Ok8pw6 = (Na0iu6 & Ql8pw6);
assign Ql8pw6 = (~(Rs4ju6 & vis_r8_o[15]));
assign Na0iu6 = (Xl8pw6 & Em8pw6);
assign Em8pw6 = (Lm8pw6 & Sm8pw6);
assign Sm8pw6 = (Zm8pw6 & Gn8pw6);
assign Gn8pw6 = (~(V6now6 & vis_r2_o[15]));
assign Zm8pw6 = (~(C7now6 & vis_r6_o[15]));
assign Lm8pw6 = (Nn8pw6 & Un8pw6);
assign Un8pw6 = (~(X7now6 & vis_r5_o[15]));
assign Nn8pw6 = (~(E8now6 & vis_r4_o[15]));
assign Xl8pw6 = (Bo8pw6 & Io8pw6);
assign Io8pw6 = (Po8pw6 & Wo8pw6);
assign Wo8pw6 = (~(N9now6 & vis_r1_o[15]));
assign Po8pw6 = (~(U9now6 & vis_r0_o[15]));
assign Bo8pw6 = (Dp8pw6 & Kp8pw6);
assign Kp8pw6 = (~(Panow6 & vis_r3_o[15]));
assign Dp8pw6 = (~(Wanow6 & vis_r7_o[15]));
assign Sfmiu6 = (!Fkfpw6[15]);
assign Bh8pw6 = (~(Eafpw6[15] & A3iiu6));
assign HADDR[14] = (Ze9iu6 ? Tugpw6[12] : Jshpw6[14]);
assign Tugpw6[12] = (~(Rp8pw6 & Yp8pw6));
assign Yp8pw6 = (~(N5fpw6[13] & Sdaiu6));
assign Rp8pw6 = (Fq8pw6 & Mq8pw6);
assign Mq8pw6 = (T2iiu6 | Xm0iu6);
assign Xm0iu6 = (Mm4ju6 ? Tq8pw6 : Kimiu6);
assign Tq8pw6 = (Ar8pw6 & Hr8pw6);
assign Hr8pw6 = (Or8pw6 & Vr8pw6);
assign Vr8pw6 = (Cs8pw6 & Js8pw6);
assign Js8pw6 = (~(Jo4ju6 & vis_r14_o[14]));
assign Cs8pw6 = (Qs8pw6 & Xs8pw6);
assign Xs8pw6 = (~(Ep4ju6 & vis_psp_o[12]));
assign Qs8pw6 = (~(Lp4ju6 & vis_msp_o[12]));
assign Or8pw6 = (Et8pw6 & Lt8pw6);
assign Lt8pw6 = (~(Gq4ju6 & vis_r12_o[14]));
assign Et8pw6 = (~(Nq4ju6 & vis_r11_o[14]));
assign Ar8pw6 = (St8pw6 & Zt8pw6);
assign Zt8pw6 = (Gu8pw6 & Nu8pw6);
assign Nu8pw6 = (~(Wr4ju6 & vis_r10_o[14]));
assign Gu8pw6 = (~(Ds4ju6 & vis_r9_o[14]));
assign St8pw6 = (Ua0iu6 & Uu8pw6);
assign Uu8pw6 = (~(Rs4ju6 & vis_r8_o[14]));
assign Ua0iu6 = (Bv8pw6 & Iv8pw6);
assign Iv8pw6 = (Pv8pw6 & Wv8pw6);
assign Wv8pw6 = (Dw8pw6 & Kw8pw6);
assign Kw8pw6 = (~(V6now6 & vis_r2_o[14]));
assign Dw8pw6 = (~(C7now6 & vis_r6_o[14]));
assign Pv8pw6 = (Rw8pw6 & Yw8pw6);
assign Yw8pw6 = (~(X7now6 & vis_r5_o[14]));
assign Rw8pw6 = (~(E8now6 & vis_r4_o[14]));
assign Bv8pw6 = (Fx8pw6 & Mx8pw6);
assign Mx8pw6 = (Tx8pw6 & Ay8pw6);
assign Ay8pw6 = (~(N9now6 & vis_r1_o[14]));
assign Tx8pw6 = (~(U9now6 & vis_r0_o[14]));
assign Fx8pw6 = (Hy8pw6 & Oy8pw6);
assign Oy8pw6 = (~(Panow6 & vis_r3_o[14]));
assign Hy8pw6 = (~(Wanow6 & vis_r7_o[14]));
assign Kimiu6 = (!Fkfpw6[14]);
assign Fq8pw6 = (~(Eafpw6[14] & A3iiu6));
assign HADDR[13] = (Ze9iu6 ? Tugpw6[11] : Jshpw6[13]);
assign Tugpw6[11] = (~(Vy8pw6 & Cz8pw6));
assign Cz8pw6 = (~(N5fpw6[12] & Sdaiu6));
assign Vy8pw6 = (Jz8pw6 & Qz8pw6);
assign Qz8pw6 = (T2iiu6 | En0iu6);
assign En0iu6 = (Mm4ju6 ? Xz8pw6 : Clmiu6);
assign Xz8pw6 = (E09pw6 & L09pw6);
assign L09pw6 = (S09pw6 & Z09pw6);
assign Z09pw6 = (G19pw6 & N19pw6);
assign N19pw6 = (~(Jo4ju6 & vis_r14_o[13]));
assign G19pw6 = (U19pw6 & B29pw6);
assign B29pw6 = (~(Ep4ju6 & vis_psp_o[11]));
assign U19pw6 = (~(Lp4ju6 & vis_msp_o[11]));
assign S09pw6 = (I29pw6 & P29pw6);
assign P29pw6 = (~(Gq4ju6 & vis_r12_o[13]));
assign I29pw6 = (~(Nq4ju6 & vis_r11_o[13]));
assign E09pw6 = (W29pw6 & D39pw6);
assign D39pw6 = (K39pw6 & R39pw6);
assign R39pw6 = (~(Wr4ju6 & vis_r10_o[13]));
assign K39pw6 = (~(Ds4ju6 & vis_r9_o[13]));
assign W29pw6 = (Bb0iu6 & Y39pw6);
assign Y39pw6 = (~(Rs4ju6 & vis_r8_o[13]));
assign Bb0iu6 = (F49pw6 & M49pw6);
assign M49pw6 = (T49pw6 & A59pw6);
assign A59pw6 = (H59pw6 & O59pw6);
assign O59pw6 = (~(V6now6 & vis_r2_o[13]));
assign H59pw6 = (~(C7now6 & vis_r6_o[13]));
assign T49pw6 = (V59pw6 & C69pw6);
assign C69pw6 = (~(X7now6 & vis_r5_o[13]));
assign V59pw6 = (~(E8now6 & vis_r4_o[13]));
assign F49pw6 = (J69pw6 & Q69pw6);
assign Q69pw6 = (X69pw6 & E79pw6);
assign E79pw6 = (~(N9now6 & vis_r1_o[13]));
assign X69pw6 = (~(U9now6 & vis_r0_o[13]));
assign J69pw6 = (L79pw6 & S79pw6);
assign S79pw6 = (~(Panow6 & vis_r3_o[13]));
assign L79pw6 = (~(Wanow6 & vis_r7_o[13]));
assign Clmiu6 = (!Fkfpw6[13]);
assign Jz8pw6 = (~(Eafpw6[13] & A3iiu6));
assign HADDR[12] = (Ze9iu6 ? Ixdpw6 : Jshpw6[12]);
assign Ixdpw6 = (~(Z79pw6 & G89pw6));
assign G89pw6 = (T2iiu6 | Ln0iu6);
assign Ln0iu6 = (Cn5ju6 ? Unmiu6 : N89pw6);
assign Cn5ju6 = (!Mm4ju6);
assign Unmiu6 = (!Fkfpw6[12]);
assign N89pw6 = (U89pw6 & B99pw6);
assign B99pw6 = (I99pw6 & P99pw6);
assign P99pw6 = (W99pw6 & Da9pw6);
assign Da9pw6 = (~(Jo4ju6 & vis_r14_o[12]));
assign W99pw6 = (Ka9pw6 & Ra9pw6);
assign Ra9pw6 = (~(Ep4ju6 & vis_psp_o[10]));
assign Ep4ju6 = (Ya9pw6 & Fb9pw6);
assign Ya9pw6 = (~(Mb9pw6 | Vq2pw6));
assign Vq2pw6 = (!Vrfhu6);
assign Ka9pw6 = (~(Lp4ju6 & vis_msp_o[10]));
assign Lp4ju6 = (Tb9pw6 & Fb9pw6);
assign Tb9pw6 = (~(Mb9pw6 | Vrfhu6));
assign I99pw6 = (Ac9pw6 & Hc9pw6);
assign Hc9pw6 = (~(Gq4ju6 & vis_r12_o[12]));
assign Ac9pw6 = (~(Nq4ju6 & vis_r11_o[12]));
assign U89pw6 = (Oc9pw6 & Vc9pw6);
assign Vc9pw6 = (Cd9pw6 & Jd9pw6);
assign Jd9pw6 = (~(Wr4ju6 & vis_r10_o[12]));
assign Cd9pw6 = (~(Ds4ju6 & vis_r9_o[12]));
assign Oc9pw6 = (Ib0iu6 & Qd9pw6);
assign Qd9pw6 = (~(Rs4ju6 & vis_r8_o[12]));
assign Ib0iu6 = (Xd9pw6 & Ee9pw6);
assign Ee9pw6 = (Le9pw6 & Se9pw6);
assign Se9pw6 = (Ze9pw6 & Gf9pw6);
assign Gf9pw6 = (~(V6now6 & vis_r2_o[12]));
assign Ze9pw6 = (~(C7now6 & vis_r6_o[12]));
assign Le9pw6 = (Nf9pw6 & Uf9pw6);
assign Uf9pw6 = (~(X7now6 & vis_r5_o[12]));
assign Nf9pw6 = (~(E8now6 & vis_r4_o[12]));
assign Xd9pw6 = (Bg9pw6 & Ig9pw6);
assign Ig9pw6 = (Pg9pw6 & Wg9pw6);
assign Wg9pw6 = (~(N9now6 & vis_r1_o[12]));
assign Pg9pw6 = (~(U9now6 & vis_r0_o[12]));
assign Bg9pw6 = (Dh9pw6 & Kh9pw6);
assign Kh9pw6 = (~(Panow6 & vis_r3_o[12]));
assign Dh9pw6 = (~(Wanow6 & vis_r7_o[12]));
assign T2iiu6 = (!B7iiu6);
assign Z79pw6 = (Rh9pw6 & Yh9pw6);
assign Yh9pw6 = (~(N5fpw6[11] & Sdaiu6));
assign Rh9pw6 = (~(Eafpw6[12] & A3iiu6));
assign HADDR[0] = (~(Fi9pw6 & Mi9pw6));
assign Mi9pw6 = (~(Ti9pw6 & E4yhu6));
assign E4yhu6 = (~(Aphpw6[1] | Aphpw6[2]));
assign Ti9pw6 = (Ne3pw6 & Tnhpw6[0]);
assign Ne3pw6 = (~(Ze9iu6 | Wqzhu6));
assign Wqzhu6 = (Ho4iu6 & H9xiu6);
assign H9xiu6 = (!Eq4iu6);
assign Eq4iu6 = (Cjhpw6[3] & Iqzhu6);
assign Ho4iu6 = (Cjhpw6[2] & Iqzhu6);
assign Iqzhu6 = (Lznhu6 ^ Dtnhu6);
assign Fi9pw6 = (~(My0iu6 & Ze9iu6));
assign Ze9iu6 = (~(Aj9pw6 & Krzhu6));
assign Krzhu6 = (~(Gpzhu6 | Sqhpw6[1]));
assign Gpzhu6 = (!Sqhpw6[0]);
assign Aj9pw6 = (HMASTER & Ebxiu6);
assign Ebxiu6 = (!Jzmhu6);
assign HMASTER = (~(Ympiu6 | S18iu6));
assign S18iu6 = (Hj9pw6 & Oj9pw6);
assign Oj9pw6 = (~(Sdaiu6 | Vj9pw6));
assign Sdaiu6 = (!Ck9pw6);
assign Hj9pw6 = (Lrhiu6 & I1aiu6);
assign My0iu6 = (Jk9pw6 & J71iu6);
assign J71iu6 = (~(X71iu6 | Mnxow6));
assign Mnxow6 = (Ed3pw6 & Qk9pw6);
assign Qk9pw6 = (~(Xk9pw6 & El9pw6));
assign El9pw6 = (~(Frziu6 & Xe8iu6));
assign Xk9pw6 = (~(Es1ju6 | Vjhow6));
assign Ed3pw6 = (!X71iu6);
assign X71iu6 = (~(Ll9pw6 & Sl9pw6));
assign Sl9pw6 = (Zl9pw6 & Gm9pw6);
assign Zl9pw6 = (Mzlow6 | Nlaiu6);
assign Mzlow6 = (Ey2ju6 | Tfjiu6);
assign Ey2ju6 = (!Fd0iu6);
assign Ll9pw6 = (Nm9pw6 & He6ju6);
assign He6ju6 = (!Ww8ow6);
assign Ww8ow6 = (Tr0iu6 & Nlaiu6);
assign Nm9pw6 = (~(H3aju6 & Sq3ju6));
assign Jk9pw6 = (~(Ympiu6 | Ta3pw6));
assign Ta3pw6 = (!Ay8iu6);
assign Ay8iu6 = (~(Um9pw6 & Bn9pw6));
assign Bn9pw6 = (~(B7iiu6 & Go0iu6));
assign Go0iu6 = (Mm4ju6 ? In9pw6 : Fkfpw6[0]);
assign Mm4ju6 = (Pn9pw6 & Wn9pw6);
assign Wn9pw6 = (Do9pw6 & Ko9pw6);
assign Ko9pw6 = (Ro9pw6 & Kgaiu6);
assign Ro9pw6 = (Yo9pw6 | Fp9pw6);
assign Do9pw6 = (Mp9pw6 & Ty8ow6);
assign Ty8ow6 = (Qxaiu6 | K9aiu6);
assign Mp9pw6 = (~(Tp9pw6 & Toaiu6));
assign Toaiu6 = (Pugiu6 & Ii0iu6);
assign Tp9pw6 = (~(Nlaiu6 | Cyfpw6[4]));
assign Pn9pw6 = (Aq9pw6 & Hq9pw6);
assign Hq9pw6 = (~(Tr0iu6 & Oq9pw6));
assign Oq9pw6 = (W8aiu6 | Oiaiu6);
assign Aq9pw6 = (Vq9pw6 & Cr9pw6);
assign Cr9pw6 = (~(Jr9pw6 & Frziu6));
assign Jr9pw6 = (~(Lkaiu6 | C0ehu6));
assign Vq9pw6 = (~(Qr9pw6 & Fhaiu6));
assign Fhaiu6 = (Nlaiu6 & Mr0iu6);
assign Qr9pw6 = (~(As0iu6 | Cyfpw6[3]));
assign In9pw6 = (~(Xr9pw6 & Es9pw6));
assign Es9pw6 = (Ls9pw6 & Ss9pw6);
assign Ss9pw6 = (Zs9pw6 & Gt9pw6);
assign Gt9pw6 = (~(Jo4ju6 & vis_r14_o[0]));
assign Jo4ju6 = (~(Yo9pw6 | Nt9pw6));
assign Zs9pw6 = (~(Gq4ju6 & vis_r12_o[0]));
assign Gq4ju6 = (~(Yo9pw6 | Ut9pw6));
assign Yo9pw6 = (!Fb9pw6);
assign Fb9pw6 = (~(Ssniu6 | Fpniu6));
assign Ls9pw6 = (Bu9pw6 & Iu9pw6);
assign Iu9pw6 = (~(Nq4ju6 & vis_r11_o[0]));
assign Nq4ju6 = (~(Pu9pw6 | Fp9pw6));
assign Bu9pw6 = (~(Wr4ju6 & vis_r10_o[0]));
assign Wr4ju6 = (~(Pu9pw6 | Nt9pw6));
assign Xr9pw6 = (Wu9pw6 & Dc0iu6);
assign Dc0iu6 = (Dv9pw6 & Kv9pw6);
assign Kv9pw6 = (Rv9pw6 & Yv9pw6);
assign Yv9pw6 = (Fw9pw6 & Mw9pw6);
assign Mw9pw6 = (~(V6now6 & vis_r2_o[0]));
assign V6now6 = (~(Tw9pw6 | Nt9pw6));
assign Fw9pw6 = (~(C7now6 & vis_r6_o[0]));
assign C7now6 = (~(Ax9pw6 | Nt9pw6));
assign Nt9pw6 = (Mxuow6 | H2fpw6[0]);
assign Rv9pw6 = (Hx9pw6 & Ox9pw6);
assign Ox9pw6 = (~(X7now6 & vis_r5_o[0]));
assign X7now6 = (~(Mb9pw6 | Ax9pw6));
assign Hx9pw6 = (~(E8now6 & vis_r4_o[0]));
assign E8now6 = (~(Ut9pw6 | Ax9pw6));
assign Dv9pw6 = (Vx9pw6 & Cy9pw6);
assign Cy9pw6 = (Jy9pw6 & Qy9pw6);
assign Qy9pw6 = (~(N9now6 & vis_r1_o[0]));
assign N9now6 = (~(Mb9pw6 | Tw9pw6));
assign Jy9pw6 = (~(U9now6 & vis_r0_o[0]));
assign U9now6 = (~(Ut9pw6 | Tw9pw6));
assign Vx9pw6 = (Xy9pw6 & Ez9pw6);
assign Ez9pw6 = (~(Panow6 & vis_r3_o[0]));
assign Panow6 = (~(Fp9pw6 | Tw9pw6));
assign Tw9pw6 = (H2fpw6[2] | H2fpw6[3]);
assign Xy9pw6 = (~(Wanow6 & vis_r7_o[0]));
assign Wanow6 = (~(Fp9pw6 | Ax9pw6));
assign Ax9pw6 = (Fpniu6 | H2fpw6[3]);
assign Fpniu6 = (!H2fpw6[2]);
assign Fp9pw6 = (Vqniu6 | Mxuow6);
assign Mxuow6 = (!H2fpw6[1]);
assign Wu9pw6 = (Lz9pw6 & Sz9pw6);
assign Sz9pw6 = (~(Ds4ju6 & vis_r9_o[0]));
assign Ds4ju6 = (~(Pu9pw6 | Mb9pw6));
assign Mb9pw6 = (Vqniu6 | H2fpw6[1]);
assign Vqniu6 = (!H2fpw6[0]);
assign Lz9pw6 = (~(Rs4ju6 & vis_r8_o[0]));
assign Rs4ju6 = (~(Pu9pw6 | Ut9pw6));
assign Ut9pw6 = (H2fpw6[0] | H2fpw6[1]);
assign Pu9pw6 = (Ssniu6 | H2fpw6[2]);
assign Ssniu6 = (!H2fpw6[3]);
assign B7iiu6 = (Zz9pw6 & Ck9pw6);
assign Zz9pw6 = (~(G0apw6 & N0apw6));
assign N0apw6 = (U0apw6 & B1apw6);
assign B1apw6 = (~(Vxniu6 & Cyfpw6[0]));
assign Vxniu6 = (~(Mjfiu6 | Tr0iu6));
assign U0apw6 = (I1apw6 & P1apw6);
assign P1apw6 = (~(W1apw6 & Fq8iu6));
assign Fq8iu6 = (H4ghu6 & Nlaiu6);
assign W1apw6 = (~(Cyfpw6[3] | Y7ghu6));
assign I1apw6 = (~(F9aju6 & Kr7ow6));
assign F9aju6 = (Cyfpw6[1] & Ii0iu6);
assign G0apw6 = (D2apw6 & K2apw6);
assign K2apw6 = (Uvziu6 | Cyfpw6[5]);
assign D2apw6 = (R2apw6 & Y2apw6);
assign Y2apw6 = (~(Z6aiu6 & Y2oiu6));
assign R2apw6 = (~(F3aiu6 & Tr0iu6));
assign Um9pw6 = (~(Eafpw6[0] & A3iiu6));
assign A3iiu6 = (F3apw6 & Ck9pw6);
assign Ck9pw6 = (~(M3apw6 & T3apw6));
assign T3apw6 = (A4apw6 & H4apw6);
assign H4apw6 = (O4apw6 & V4apw6);
assign V4apw6 = (~(C5apw6 & Mfjiu6));
assign C5apw6 = (~(Sbghu6 | Cyfpw6[6]));
assign O4apw6 = (J5apw6 & Td0iu6);
assign J5apw6 = (~(Cyfpw6[7] & Q5apw6));
assign Q5apw6 = (X5apw6 | I82ju6);
assign I82ju6 = (Apaiu6 & L45iu6);
assign X5apw6 = (Cyfpw6[4] ? Z6aiu6 : N1aow6);
assign N1aow6 = (Wwziu6 & Sijiu6);
assign Sijiu6 = (!N2ghu6);
assign A4apw6 = (E6apw6 & L6apw6);
assign L6apw6 = (~(S6apw6 & Gwyiu6));
assign S6apw6 = (~(Kq0iu6 | Ae0iu6));
assign E6apw6 = (Z6apw6 & G7apw6);
assign G7apw6 = (~(N7apw6 & Hzziu6));
assign N7apw6 = (~(Tr0iu6 | H4ghu6));
assign Z6apw6 = (~(U7apw6 & B8apw6));
assign U7apw6 = (~(Nloiu6 | Cyfpw6[4]));
assign M3apw6 = (I8apw6 & P8apw6);
assign P8apw6 = (W8apw6 & Cq3pw6);
assign Cq3pw6 = (Mjfiu6 | Mr0iu6);
assign Mjfiu6 = (!Xzmiu6);
assign Xzmiu6 = (Ii0iu6 & Tfjiu6);
assign W8apw6 = (D9apw6 & Oq1ju6);
assign Oq1ju6 = (~(Qe8iu6 & G47ow6));
assign G47ow6 = (Xe8iu6 & Tfjiu6);
assign Qe8iu6 = (~(P1bow6 | C0ehu6));
assign D9apw6 = (~(K9apw6 & R9apw6));
assign R9apw6 = (~(Qxaiu6 | Cyfpw6[5]));
assign K9apw6 = (Yljiu6 & Qyniu6);
assign I8apw6 = (Y9apw6 & Rcziu6);
assign Rcziu6 = (Faapw6 & Oe8ow6);
assign Oe8ow6 = (K9aiu6 | Tr0iu6);
assign Faapw6 = (~(Gwyiu6 & Maapw6));
assign Maapw6 = (Vbiow6 | Y0jiu6);
assign Y0jiu6 = (H4ghu6 & It2ju6);
assign Vbiow6 = (~(Xojiu6 | Kq0iu6));
assign Y9apw6 = (Taapw6 & Abapw6);
assign Abapw6 = (~(Hbapw6 & Hiaiu6));
assign Hbapw6 = (~(Iuniu6 | Nlaiu6));
assign Taapw6 = (~(Ls1ju6 & Md0iu6));
assign Md0iu6 = (~(Cyfpw6[0] | Cyfpw6[4]));
assign Ls1ju6 = (Apaiu6 & Jjhiu6);
assign Apaiu6 = (~(Jcaiu6 | Sbghu6));
assign F3apw6 = (~(Obapw6 & Vbapw6));
assign Vbapw6 = (Ccapw6 & Jcapw6);
assign Jcapw6 = (~(Jf6ju6 | Pthiu6));
assign Jf6ju6 = (Tr0iu6 & Ii0iu6);
assign Ccapw6 = (Qcapw6 & Xcapw6);
assign Xcapw6 = (~(Edapw6 & Owoiu6));
assign Owoiu6 = (Cyfpw6[3] & Xe8iu6);
assign Edapw6 = (~(Cyfpw6[4] | Y7ghu6));
assign Qcapw6 = (~(H4ghu6 & Ldapw6));
assign Ldapw6 = (Cyfpw6[4] | A3aju6);
assign A3aju6 = (Cyfpw6[0] & Cyfpw6[1]);
assign Obapw6 = (Sdapw6 & Zdapw6);
assign Zdapw6 = (Geapw6 & Wh7ju6);
assign Wh7ju6 = (O60ju6 | Cyfpw6[0]);
assign O60ju6 = (!Vjhow6);
assign Vjhow6 = (H4ghu6 & Cyfpw6[5]);
assign Geapw6 = (Tfjiu6 | Lkaiu6);
assign Sdapw6 = (Cyfpw6[7] & Neapw6);
assign Neapw6 = (Qxaiu6 | Tr0iu6);
assign Ympiu6 = (!Ob3pw6);
assign Ob3pw6 = (~(Ueapw6 & Bfapw6));
assign Bfapw6 = (Aphiu6 & Ifapw6);
assign Ifapw6 = (~(Pfapw6 & Srhiu6));
assign Srhiu6 = (~(B7qow6 & Et8iu6));
assign Pfapw6 = (vis_pc_o[0] ? Dgapw6 : Wfapw6);
assign Dgapw6 = (Kgapw6 & Rgapw6);
assign Rgapw6 = (~(Juzhu6 & Ophiu6));
assign Juzhu6 = (~(Sufpw6[1] & Ygapw6));
assign Kgapw6 = (Jjhiu6 | Dxfhu6);
assign Wfapw6 = (~(Ophiu6 & N6piu6));
assign N6piu6 = (!Pkciu6);
assign Pkciu6 = (Sufpw6[0] & Ygapw6);
assign Ophiu6 = (~(B7qow6 & U6qow6));
assign U6qow6 = (!Gu8iu6);
assign Gu8iu6 = (Kgaiu6 & Fhapw6);
assign Fhapw6 = (~(Yp8iu6 & Hzziu6));
assign Yp8iu6 = (Cyfpw6[5] & Nlaiu6);
assign Kgaiu6 = (!Uoziu6);
assign Uoziu6 = (L78ju6 & Y7ghu6);
assign Aphiu6 = (I1aiu6 & Dp8iu6);
assign Dp8iu6 = (!LOCKUP);
assign LOCKUP = (~(Mhapw6 & Thapw6));
assign Thapw6 = (~(Aiapw6 & H3aju6));
assign Aiapw6 = (Mfjiu6 & Sbghu6);
assign Mhapw6 = (Hiapw6 & Oiapw6);
assign Oiapw6 = (~(Omyiu6 & Viapw6));
assign Viapw6 = (~(Cjapw6 & Jjapw6));
assign Jjapw6 = (~(Qjapw6 & Xjapw6));
assign Xjapw6 = (Kxziu6 & Kr7ow6);
assign Kr7ow6 = (~(Vwaiu6 | H4ghu6));
assign Qjapw6 = (~(Ruaiu6 | Wfoiu6));
assign Ruaiu6 = (!V9ghu6);
assign Cjapw6 = (~(Ekapw6 & Lkapw6));
assign Lkapw6 = (~(Y7ghu6 | H4ghu6));
assign Ekapw6 = (~(Qjaiu6 | Cyfpw6[5]));
assign Hiapw6 = (~(V9ghu6 & Skapw6));
assign Skapw6 = (~(Xxaiu6 & Zkapw6));
assign Xxaiu6 = (Glapw6 & Nlapw6);
assign Nlapw6 = (Ulapw6 & Bmapw6);
assign Bmapw6 = (~(Imapw6 & Buaow6));
assign Imapw6 = (~(Ntgiu6 | P0biu6));
assign P0biu6 = (Pmapw6 & Wmapw6);
assign Wmapw6 = (~(Dnapw6 & Knapw6));
assign Knapw6 = (Sbrow6 | B3gpw6[1]);
assign Dnapw6 = (Rnapw6 & Gcrow6);
assign Gcrow6 = (~(Ynapw6 & Foapw6));
assign Foapw6 = (Moapw6 & Toapw6);
assign Toapw6 = (Apapw6 & Hpapw6);
assign Hpapw6 = (Opapw6 & Vpapw6);
assign Vpapw6 = (Cqapw6 & Oyfiu6);
assign Cqapw6 = (~(Arfiu6 | Ahbiu6));
assign Opapw6 = (~(Lhdiu6 | Nbdiu6));
assign Apapw6 = (Jqapw6 & Qqapw6);
assign Qqapw6 = (~(Jndiu6 | Kkdiu6));
assign Jqapw6 = (~(V5giu6 | Iqdiu6));
assign Moapw6 = (Xqapw6 & Erapw6);
assign Erapw6 = (Lrapw6 & Srapw6);
assign Srapw6 = (Zrapw6 & Coxiu6);
assign Zrapw6 = (~(Bggiu6 | Z7giu6));
assign Lrapw6 = (~(Umgiu6 | Odfiu6));
assign Xqapw6 = (Gsapw6 & Nsapw6);
assign Nsapw6 = (~(Hl7iu6 | Yogiu6));
assign Gsapw6 = (~(Ajgiu6 | Qrgiu6));
assign Ynapw6 = (Usapw6 & Btapw6);
assign Btapw6 = (Itapw6 & Ptapw6);
assign Ptapw6 = (Wtapw6 & Duapw6);
assign Duapw6 = (Kuapw6 & Giyiu6);
assign Kuapw6 = (~(Webiu6 | Rhgiu6));
assign Wtapw6 = (~(Ivfiu6 | Etfiu6));
assign Ivfiu6 = (!Ubyiu6);
assign Itapw6 = (Ruapw6 & Yuapw6);
assign Yuapw6 = (~(O8diu6 | Mxfiu6));
assign Ruapw6 = (~(N1giu6 | Mediu6));
assign Usapw6 = (Fvapw6 & Mvapw6);
assign Mvapw6 = (Tvapw6 & Awapw6);
assign Awapw6 = (~(R3giu6 | Hwhiu6));
assign Tvapw6 = (~(Hcgiu6 | Dagiu6));
assign Hcgiu6 = (!Spxiu6);
assign Fvapw6 = (Hwapw6 & Owapw6);
assign Owapw6 = (~(G9fiu6 | Eegiu6));
assign Hwapw6 = (~(Sffiu6 | Kbfiu6));
assign Rnapw6 = (~(Vwapw6 & Cxapw6));
assign Cxapw6 = (~(Sbrow6 & B3gpw6[1]));
assign Sbrow6 = (Jxapw6 & Qxapw6);
assign Qxapw6 = (Xxapw6 & Eyapw6);
assign Eyapw6 = (Lyapw6 & Syapw6);
assign Syapw6 = (Zyapw6 & Gzapw6);
assign Gzapw6 = (Nzapw6 & Uzapw6);
assign Uzapw6 = (~(B3gpw6[1] & Qrgiu6));
assign Nzapw6 = (B0bpw6 & I0bpw6);
assign I0bpw6 = (~(L1gpw6[1] & Rhgiu6));
assign B0bpw6 = (~(H8gpw6[1] & Ajgiu6));
assign Zyapw6 = (P0bpw6 & W0bpw6);
assign W0bpw6 = (U2uow6 | Ucxiu6);
assign U2uow6 = (!R4gpw6[1]);
assign P0bpw6 = (~(R4gpw6[3] & Yogiu6));
assign Lyapw6 = (D1bpw6 & K1bpw6);
assign K1bpw6 = (R1bpw6 & Y1bpw6);
assign Y1bpw6 = (Fytow6 | Agxiu6);
assign Fytow6 = (!R4gpw6[5]);
assign R1bpw6 = (Yxtow6 | Qhxiu6);
assign Qhxiu6 = (!Sffiu6);
assign Yxtow6 = (!R4gpw6[7]);
assign D1bpw6 = (F2bpw6 & M2bpw6);
assign M2bpw6 = (~(R4gpw6[9] & Odfiu6));
assign F2bpw6 = (Yqtow6 | Wkxiu6);
assign Wkxiu6 = (!Kbfiu6);
assign Yqtow6 = (!R4gpw6[11]);
assign Xxapw6 = (T2bpw6 & A3bpw6);
assign A3bpw6 = (H3bpw6 & O3bpw6);
assign O3bpw6 = (V3bpw6 & C4bpw6);
assign C4bpw6 = (Mrtow6 | Mmxiu6);
assign Mmxiu6 = (!G9fiu6);
assign Mrtow6 = (!R4gpw6[13]);
assign V3bpw6 = (J4bpw6 & Q4bpw6);
assign Q4bpw6 = (Frtow6 | Coxiu6);
assign Frtow6 = (!R4gpw6[15]);
assign J4bpw6 = (Xluow6 | Gfgiu6);
assign Xluow6 = (!R4gpw6[17]);
assign H3bpw6 = (X4bpw6 & E5bpw6);
assign E5bpw6 = (Qluow6 | Jdgiu6);
assign Qluow6 = (!R4gpw6[19]);
assign X4bpw6 = (Pouow6 | Spxiu6);
assign Pouow6 = (!R4gpw6[21]);
assign T2bpw6 = (L5bpw6 & S5bpw6);
assign S5bpw6 = (Z5bpw6 & G6bpw6);
assign G6bpw6 = (Wouow6 | Irxiu6);
assign Wouow6 = (!R4gpw6[23]);
assign Z5bpw6 = (~(R4gpw6[25] & Z7giu6));
assign L5bpw6 = (N6bpw6 & U6bpw6);
assign U6bpw6 = (Ihuow6 | Ouxiu6);
assign Ihuow6 = (!R4gpw6[27]);
assign N6bpw6 = (~(R4gpw6[29] & R3giu6));
assign Jxapw6 = (B7bpw6 & I7bpw6);
assign I7bpw6 = (P7bpw6 & W7bpw6);
assign W7bpw6 = (D8bpw6 & K8bpw6);
assign K8bpw6 = (R8bpw6 & Y8bpw6);
assign Y8bpw6 = (Mcuow6 | Nxxiu6);
assign Mcuow6 = (!R4gpw6[31]);
assign R8bpw6 = (F9bpw6 & M9bpw6);
assign M9bpw6 = (~(R4gpw6[33] & Hwhiu6));
assign F9bpw6 = (Dksow6 | M0yiu6);
assign M0yiu6 = (!Iqdiu6);
assign Dksow6 = (!R4gpw6[35]);
assign D8bpw6 = (T9bpw6 & Aabpw6);
assign Aabpw6 = (Ehsow6 | C2yiu6);
assign C2yiu6 = (!Jndiu6);
assign Ehsow6 = (!R4gpw6[37]);
assign T9bpw6 = (~(R4gpw6[39] & Kkdiu6));
assign P7bpw6 = (Habpw6 & Oabpw6);
assign Oabpw6 = (Vabpw6 & Cbbpw6);
assign Cbbpw6 = (~(R4gpw6[41] & Lhdiu6));
assign Vabpw6 = (Q9sow6 | Y6yiu6);
assign Y6yiu6 = (!Mediu6);
assign Q9sow6 = (!R4gpw6[43]);
assign Habpw6 = (Jbbpw6 & Qbbpw6);
assign Qbbpw6 = (Ubsow6 | O8yiu6);
assign O8yiu6 = (!Nbdiu6);
assign Ubsow6 = (!R4gpw6[45]);
assign Jbbpw6 = (~(R4gpw6[47] & O8diu6));
assign B7bpw6 = (Xbbpw6 & Ecbpw6);
assign Ecbpw6 = (Lcbpw6 & Scbpw6);
assign Scbpw6 = (Zcbpw6 & Gdbpw6);
assign Gdbpw6 = (Otsow6 | Oyfiu6);
assign Otsow6 = (!R4gpw6[49]);
assign Zcbpw6 = (Htsow6 | Rwfiu6);
assign Htsow6 = (!R4gpw6[51]);
assign Lcbpw6 = (Ndbpw6 & Udbpw6);
assign Udbpw6 = (Vtsow6 | Ubyiu6);
assign Vtsow6 = (!R4gpw6[53]);
assign Ndbpw6 = (Cusow6 | Kdyiu6);
assign Cusow6 = (!R4gpw6[55]);
assign Xbbpw6 = (Bebpw6 & Iebpw6);
assign Iebpw6 = (Pebpw6 & Webpw6);
assign Webpw6 = (~(R4gpw6[57] & Arfiu6));
assign Pebpw6 = (V7tow6 | Qgyiu6);
assign V7tow6 = (!R4gpw6[59]);
assign Bebpw6 = (Dfbpw6 & Kfbpw6);
assign Kfbpw6 = (E2tow6 | Giyiu6);
assign Giyiu6 = (!Lyhiu6);
assign E2tow6 = (!R4gpw6[61]);
assign Dfbpw6 = (~(R4gpw6[63] & Webiu6));
assign Vwapw6 = (Idrow6 & Xglow6);
assign Xglow6 = (!B3gpw6[0]);
assign Idrow6 = (~(Rfbpw6 & Yfbpw6));
assign Yfbpw6 = (Fgbpw6 & Mgbpw6);
assign Mgbpw6 = (Tgbpw6 & Ahbpw6);
assign Ahbpw6 = (Hhbpw6 & Ohbpw6);
assign Ohbpw6 = (Vhbpw6 & Cibpw6);
assign Cibpw6 = (~(B3gpw6[0] & Qrgiu6));
assign Qrgiu6 = (F8row6 & Jibpw6);
assign Vhbpw6 = (Qibpw6 & Xibpw6);
assign Xibpw6 = (~(L1gpw6[0] & Rhgiu6));
assign Rhgiu6 = (Ejbpw6 & A9row6);
assign Ejbpw6 = (Ljbpw6 & H9row6);
assign Qibpw6 = (~(H8gpw6[0] & Ajgiu6));
assign Ajgiu6 = (F8row6 & Ljbpw6);
assign F8row6 = (Sjbpw6 & H9row6);
assign Hhbpw6 = (Zjbpw6 & Gkbpw6);
assign Gkbpw6 = (B3uow6 | Ucxiu6);
assign Ucxiu6 = (!Hl7iu6);
assign Hl7iu6 = (Nkbpw6 & Ukbpw6);
assign B3uow6 = (!R4gpw6[0]);
assign Zjbpw6 = (~(R4gpw6[2] & Yogiu6));
assign Yogiu6 = (~(Blbpw6 | Ilbpw6));
assign Tgbpw6 = (Plbpw6 & Wlbpw6);
assign Wlbpw6 = (Dmbpw6 & Kmbpw6);
assign Kmbpw6 = (J0uow6 | Agxiu6);
assign Agxiu6 = (!Umgiu6);
assign Umgiu6 = (Nkbpw6 & A9row6);
assign J0uow6 = (!R4gpw6[4]);
assign Dmbpw6 = (~(R4gpw6[6] & Sffiu6));
assign Sffiu6 = (Nkbpw6 & Sjbpw6);
assign Nkbpw6 = (!Blbpw6);
assign Blbpw6 = (~(Rmbpw6 & M8row6));
assign Plbpw6 = (Ymbpw6 & Fnbpw6);
assign Fnbpw6 = (~(R4gpw6[8] & Odfiu6));
assign Odfiu6 = (~(Mnbpw6 | Tnbpw6));
assign Ymbpw6 = (~(R4gpw6[10] & Kbfiu6));
assign Kbfiu6 = (Aobpw6 & Hobpw6);
assign Fgbpw6 = (Oobpw6 & Vobpw6);
assign Vobpw6 = (Cpbpw6 & Jpbpw6);
assign Jpbpw6 = (Qpbpw6 & Xpbpw6);
assign Xpbpw6 = (~(R4gpw6[12] & G9fiu6));
assign G9fiu6 = (~(Mnbpw6 | Eqbpw6));
assign Mnbpw6 = (!Aobpw6);
assign Qpbpw6 = (Lqbpw6 & Sqbpw6);
assign Sqbpw6 = (Qttow6 | Coxiu6);
assign Coxiu6 = (!C7fiu6);
assign C7fiu6 = (Aobpw6 & Sjbpw6);
assign Aobpw6 = (Zqbpw6 & Rmbpw6);
assign Qttow6 = (!R4gpw6[14]);
assign Lqbpw6 = (Iouow6 | Gfgiu6);
assign Gfgiu6 = (!Bggiu6);
assign Bggiu6 = (~(Grbpw6 | Tnbpw6));
assign Iouow6 = (!R4gpw6[16]);
assign Cpbpw6 = (Nrbpw6 & Urbpw6);
assign Urbpw6 = (~(R4gpw6[18] & Eegiu6));
assign Eegiu6 = (!Jdgiu6);
assign Jdgiu6 = (Grbpw6 | Ilbpw6);
assign Nrbpw6 = (Aruow6 | Spxiu6);
assign Spxiu6 = (Grbpw6 | Eqbpw6);
assign Aruow6 = (!R4gpw6[20]);
assign Oobpw6 = (Bsbpw6 & Isbpw6);
assign Isbpw6 = (Psbpw6 & Wsbpw6);
assign Wsbpw6 = (~(R4gpw6[22] & Dagiu6));
assign Dagiu6 = (!Irxiu6);
assign Irxiu6 = (Grbpw6 | Dtbpw6);
assign Grbpw6 = (~(Rmbpw6 & Jibpw6));
assign Psbpw6 = (~(R4gpw6[24] & Z7giu6));
assign Z7giu6 = (!Ysxiu6);
assign Ysxiu6 = (~(Ktbpw6 & Rmbpw6));
assign Ktbpw6 = (Ljbpw6 & Ukbpw6);
assign Bsbpw6 = (Rtbpw6 & Ytbpw6);
assign Ytbpw6 = (~(R4gpw6[26] & V5giu6));
assign V5giu6 = (!Ouxiu6);
assign Ouxiu6 = (~(Fubpw6 & Rmbpw6));
assign Fubpw6 = (Ljbpw6 & Hobpw6);
assign Rtbpw6 = (~(R4gpw6[28] & R3giu6));
assign R3giu6 = (Mubpw6 & Rmbpw6);
assign Mubpw6 = (A9row6 & Ljbpw6);
assign Rfbpw6 = (Tubpw6 & Avbpw6);
assign Avbpw6 = (Hvbpw6 & Ovbpw6);
assign Ovbpw6 = (Vvbpw6 & Cwbpw6);
assign Cwbpw6 = (Jwbpw6 & Qwbpw6);
assign Qwbpw6 = (~(R4gpw6[30] & N1giu6));
assign N1giu6 = (!Nxxiu6);
assign Nxxiu6 = (~(Xwbpw6 & Rmbpw6));
assign Rmbpw6 = (vis_ipsr_o[4] & Vhbiu6);
assign Xwbpw6 = (Sjbpw6 & Ljbpw6);
assign Jwbpw6 = (Exbpw6 & Lxbpw6);
assign Lxbpw6 = (~(R4gpw6[32] & Hwhiu6));
assign Hwhiu6 = (~(Sxbpw6 | Tnbpw6));
assign Exbpw6 = (~(R4gpw6[34] & Iqdiu6));
assign Iqdiu6 = (Zxbpw6 & Hobpw6);
assign Vvbpw6 = (Gybpw6 & Nybpw6);
assign Nybpw6 = (~(R4gpw6[36] & Jndiu6));
assign Jndiu6 = (Zxbpw6 & A9row6);
assign Gybpw6 = (Lhsow6 | S3yiu6);
assign S3yiu6 = (!Kkdiu6);
assign Kkdiu6 = (Sjbpw6 & Zxbpw6);
assign Zxbpw6 = (!Sxbpw6);
assign Sxbpw6 = (~(Uybpw6 & M8row6));
assign Lhsow6 = (!R4gpw6[38]);
assign Hvbpw6 = (Bzbpw6 & Izbpw6);
assign Izbpw6 = (Pzbpw6 & Wzbpw6);
assign Wzbpw6 = (~(R4gpw6[40] & Lhdiu6));
assign Lhdiu6 = (~(D0cpw6 | Tnbpw6));
assign Pzbpw6 = (~(R4gpw6[42] & Mediu6));
assign Mediu6 = (K0cpw6 & Hobpw6);
assign Bzbpw6 = (R0cpw6 & Y0cpw6);
assign Y0cpw6 = (~(R4gpw6[44] & Nbdiu6));
assign Nbdiu6 = (~(Eqbpw6 | D0cpw6));
assign D0cpw6 = (!K0cpw6);
assign R0cpw6 = (Bcsow6 | Eayiu6);
assign Eayiu6 = (!O8diu6);
assign O8diu6 = (Sjbpw6 & K0cpw6);
assign K0cpw6 = (Zqbpw6 & Uybpw6);
assign Zqbpw6 = (~(Tfciu6 | vis_ipsr_o[3]));
assign Bcsow6 = (!R4gpw6[46]);
assign Tubpw6 = (F1cpw6 & M1cpw6);
assign M1cpw6 = (T1cpw6 & A2cpw6);
assign A2cpw6 = (H2cpw6 & O2cpw6);
assign O2cpw6 = (Yysow6 | Oyfiu6);
assign Oyfiu6 = (!Jzfiu6);
assign Jzfiu6 = (~(V2cpw6 | Tnbpw6));
assign Tnbpw6 = (!Ukbpw6);
assign Yysow6 = (!R4gpw6[48]);
assign H2cpw6 = (~(R4gpw6[50] & Mxfiu6));
assign Mxfiu6 = (!Rwfiu6);
assign Rwfiu6 = (V2cpw6 | Ilbpw6);
assign T1cpw6 = (C3cpw6 & J3cpw6);
assign J3cpw6 = (Uwsow6 | Ubyiu6);
assign Ubyiu6 = (Eqbpw6 | V2cpw6);
assign Eqbpw6 = (!A9row6);
assign Uwsow6 = (!R4gpw6[52]);
assign C3cpw6 = (~(R4gpw6[54] & Etfiu6));
assign Etfiu6 = (!Kdyiu6);
assign Kdyiu6 = (Dtbpw6 | V2cpw6);
assign V2cpw6 = (~(Jibpw6 & Uybpw6));
assign Jibpw6 = (~(Ngfiu6 | vis_ipsr_o[2]));
assign Dtbpw6 = (!Sjbpw6);
assign F1cpw6 = (Q3cpw6 & X3cpw6);
assign X3cpw6 = (E4cpw6 & L4cpw6);
assign L4cpw6 = (~(R4gpw6[56] & Arfiu6));
assign Arfiu6 = (!Afyiu6);
assign Afyiu6 = (~(S4cpw6 & Ljbpw6));
assign S4cpw6 = (Uybpw6 & Ukbpw6);
assign E4cpw6 = (~(R4gpw6[58] & Ahbiu6));
assign Ahbiu6 = (!Qgyiu6);
assign Qgyiu6 = (~(Z4cpw6 & Ljbpw6));
assign Z4cpw6 = (Uybpw6 & Hobpw6);
assign Hobpw6 = (!Ilbpw6);
assign Ilbpw6 = (~(vis_ipsr_o[0] & Siciu6));
assign Q3cpw6 = (G5cpw6 & N5cpw6);
assign N5cpw6 = (~(R4gpw6[60] & Lyhiu6));
assign Lyhiu6 = (U5cpw6 & A9row6);
assign G5cpw6 = (~(R4gpw6[62] & Webiu6));
assign Webiu6 = (U5cpw6 & Sjbpw6);
assign U5cpw6 = (Ljbpw6 & Uybpw6);
assign Uybpw6 = (~(Vhbiu6 | vis_ipsr_o[4]));
assign Vhbiu6 = (!vis_ipsr_o[5]);
assign Ljbpw6 = (~(Ngfiu6 | Tfciu6));
assign Tfciu6 = (!vis_ipsr_o[2]);
assign Ngfiu6 = (!vis_ipsr_o[3]);
assign Pmapw6 = (~(B6cpw6 | vis_primask_o));
assign B6cpw6 = (I6cpw6 & H9row6);
assign I6cpw6 = (M8row6 & P6cpw6);
assign P6cpw6 = (A9row6 | Sjbpw6);
assign Sjbpw6 = (vis_ipsr_o[1] & vis_ipsr_o[0]);
assign A9row6 = (~(Siciu6 | vis_ipsr_o[0]));
assign Siciu6 = (!vis_ipsr_o[1]);
assign Ulapw6 = (~(W6cpw6 & D7cpw6));
assign D7cpw6 = (K7cpw6 & Kxziu6);
assign K7cpw6 = (~(R75iu6 | Hbbow6));
assign R75iu6 = (!Omyiu6);
assign W6cpw6 = (L78ju6 & Frziu6);
assign Glapw6 = (Erhiu6 & R7cpw6);
assign R7cpw6 = (~(Jxaiu6 & Y7cpw6));
assign Y7cpw6 = (~(F8cpw6 & M8cpw6));
assign M8cpw6 = (~(T8cpw6 & A9cpw6));
assign A9cpw6 = (Ftjiu6 | D7fpw6[14]);
assign T8cpw6 = (~(Xjbow6 | D7fpw6[12]));
assign Xjbow6 = (D7fpw6[14] & S1ehu6);
assign F8cpw6 = (~(Y40ju6 | Jiiiu6));
assign Jxaiu6 = (H9cpw6 & O9cpw6);
assign O9cpw6 = (~(Y2oiu6 | Jcaiu6));
assign H9cpw6 = (~(Wfoiu6 | Ccoiu6));
assign I1aiu6 = (~(Pu1ju6 & B8apw6));
assign Ueapw6 = (Erhiu6 & Lrhiu6);
assign Lrhiu6 = (V9cpw6 & Cacpw6);
assign Cacpw6 = (Jacpw6 & Qacpw6);
assign Qacpw6 = (Xacpw6 & Uloiu6);
assign Uloiu6 = (~(Ebcpw6 & N2ghu6));
assign Ebcpw6 = (Whfiu6 & D6kiu6);
assign Whfiu6 = (Cyfpw6[3] & Cyfpw6[5]);
assign Xacpw6 = (Kz6ow6 & Td0iu6);
assign Td0iu6 = (~(Omyiu6 & Pfiow6));
assign Pfiow6 = (Lbcpw6 & Oiaiu6);
assign Lbcpw6 = (Sq3ju6 & Cyfpw6[5]);
assign Kz6ow6 = (~(Sbcpw6 & Pthiu6));
assign Sbcpw6 = (~(Jojiu6 | Ii0iu6));
assign Jojiu6 = (!Pu1ju6);
assign Pu1ju6 = (~(Mr0iu6 | K9aiu6));
assign Jacpw6 = (~(Zbcpw6 | Iepiu6));
assign Iepiu6 = (W8aiu6 & Ldoiu6);
assign Zbcpw6 = (Wp0iu6 & D6kiu6);
assign V9cpw6 = (Gccpw6 & Nccpw6);
assign Nccpw6 = (Zkapw6 & Uccpw6);
assign Uccpw6 = (~(Ae0iu6 & Bdcpw6));
assign Bdcpw6 = (~(Idcpw6 & Pdcpw6));
assign Pdcpw6 = (Wdcpw6 & Decpw6);
assign Decpw6 = (~(N3ziu6 & Kecpw6));
assign Kecpw6 = (Y2oiu6 | X97ow6);
assign N3ziu6 = (Yljiu6 & Nlaiu6);
assign Wdcpw6 = (Recpw6 & Iw8ow6);
assign Iw8ow6 = (~(Yecpw6 & Wwziu6));
assign Wwziu6 = (!Nloiu6);
assign Nloiu6 = (~(D6kiu6 & H4ghu6));
assign Yecpw6 = (~(Y2oiu6 | Xe8iu6));
assign Recpw6 = (~(Ffcpw6 & Pt2ju6));
assign Ffcpw6 = (~(C0ehu6 | Cyfpw6[6]));
assign Idcpw6 = (Mfcpw6 & Tfcpw6);
assign Tfcpw6 = (Qjaiu6 | Kw0ju6);
assign Mfcpw6 = (Agcpw6 & Hgcpw6);
assign Hgcpw6 = (~(S6aiu6 & Ogcpw6));
assign Ogcpw6 = (~(Owaiu6 & Vgcpw6));
assign Vgcpw6 = (Xmliu6 | Cyfpw6[0]);
assign Owaiu6 = (!Cp3ju6);
assign Agcpw6 = (~(Chcpw6 & K9aiu6));
assign Chcpw6 = (~(Jhcpw6 & Qhcpw6));
assign Qhcpw6 = (~(L45iu6 & Oiaiu6));
assign L45iu6 = (~(Gm9pw6 | Cyfpw6[4]));
assign Gm9pw6 = (Cyfpw6[3] | C0ehu6);
assign Jhcpw6 = (Lkaiu6 | Mr0iu6);
assign Zkapw6 = (~(Xhcpw6 & Eicpw6));
assign Eicpw6 = (~(Knaiu6 | Cyfpw6[5]));
assign Xhcpw6 = (~(As0iu6 | Qxaiu6));
assign Gccpw6 = (Licpw6 & Sicpw6);
assign Sicpw6 = (~(Zicpw6 & Mmjiu6));
assign Mmjiu6 = (!Qu7ow6);
assign Qu7ow6 = (Nsaiu6 | Pxyiu6);
assign Pxyiu6 = (~(Gjcpw6 & vis_pc_o[2]));
assign Gjcpw6 = (Qqdhu6 & El1ju6);
assign Nsaiu6 = (~(Njcpw6 & Q5aiu6));
assign Njcpw6 = (El1ju6 | E6phu6);
assign El1ju6 = (!Stdhu6);
assign Zicpw6 = (~(Qjaiu6 | Kw0ju6));
assign Kw0ju6 = (~(I30ju6 & Ii0iu6));
assign I30ju6 = (~(R2aiu6 | Dxziu6));
assign Dxziu6 = (!Xojiu6);
assign Xojiu6 = (~(Ujcpw6 & Bkcpw6));
assign Bkcpw6 = (Ikcpw6 & Pkcpw6);
assign Pkcpw6 = (~(Xkhow6 | Qbiiu6));
assign Qbiiu6 = (S8fpw6[9] & S8fpw6[8]);
assign Xkhow6 = (S8fpw6[7] & L28ow6);
assign L28ow6 = (G55iu6 | S8fpw6[6]);
assign Ikcpw6 = (Wj7ow6 & G7iow6);
assign G7iow6 = (~(S8fpw6[6] & G55iu6));
assign G55iu6 = (Wkcpw6 | S8fpw6[5]);
assign Wj7ow6 = (~(S8fpw6[5] & Wkcpw6));
assign Wkcpw6 = (!Zoyiu6);
assign Zoyiu6 = (N55iu6 & Qjoiu6);
assign Ujcpw6 = (Dlcpw6 & Klcpw6);
assign Klcpw6 = (~(S8fpw6[10] & Weiiu6));
assign Dlcpw6 = (Voiiu6 & Btbow6);
assign Btbow6 = (Qjoiu6 | N55iu6);
assign N55iu6 = (~(B65iu6 | S8fpw6[11]));
assign Qjoiu6 = (!S8fpw6[4]);
assign Voiiu6 = (~(S8fpw6[11] & B65iu6));
assign B65iu6 = (Weiiu6 | S8fpw6[10]);
assign Weiiu6 = (S8fpw6[8] | S8fpw6[9]);
assign Licpw6 = (Cyfpw6[4] ? Ylcpw6 : Rlcpw6);
assign Ylcpw6 = (Ccoiu6 | Geaiu6);
assign Rlcpw6 = (Fmcpw6 & Mmcpw6);
assign Mmcpw6 = (~(Z6aiu6 & Oiaiu6));
assign Fmcpw6 = (Tmcpw6 & Ancpw6);
assign Ancpw6 = (~(Hncpw6 & K2aiu6));
assign Hncpw6 = (N2ghu6 & D6kiu6);
assign Tmcpw6 = (Jc2ju6 | R2aiu6);
assign R2aiu6 = (!W8aiu6);
assign Jc2ju6 = (!Es1ju6);
assign Es1ju6 = (Nlaiu6 & Xe8iu6);
assign GATEHCLK = (~(CDBGPWRUPACK | Oncpw6));
assign Oncpw6 = (~(E6phu6 | SLEEPING));
assign SLEEPING = (Qnghu6 & Vncpw6);
assign CODENSEQ = (~(Cocpw6 & Jocpw6));
assign Jocpw6 = (Qocpw6 & Uriiu6);
assign Qocpw6 = (~(Hrfpw6[16] | Yyfhu6));
assign Cocpw6 = (Xocpw6 & Epcpw6);
assign Epcpw6 = (~(Ppfpw6[16] & Ntfhu6));
assign Xocpw6 = (Lpcpw6 & Ygapw6);
assign Ygapw6 = (~(Spcpw6 & Gc5iu6));
assign Gc5iu6 = (!Wofiu6);
assign Wofiu6 = (~(L6aiu6 & Zpcpw6));
assign Zpcpw6 = (~(B8apw6 & D6kiu6));
assign B8apw6 = (~(Ccoiu6 | Ii0iu6));
assign Ccoiu6 = (!H3aju6);
assign H3aju6 = (Cyfpw6[7] & Xe8iu6);
assign L6aiu6 = (~(Wp0iu6 & Mfjiu6));
assign Mfjiu6 = (Cyfpw6[4] & Y7ghu6);
assign Spcpw6 = (B7qow6 & Et8iu6);
assign Et8iu6 = (U0aiu6 | Gqcpw6);
assign Gqcpw6 = (D1piu6 & Tr0iu6);
assign U0aiu6 = (Hzziu6 & Cyfpw6[0]);
assign B7qow6 = (~(Nqcpw6 & Uqcpw6));
assign Uqcpw6 = (Brcpw6 & Ircpw6);
assign Ircpw6 = (~(Prcpw6 | Nz2ju6));
assign Nz2ju6 = (F23ju6 & D31ju6);
assign D31ju6 = (Cyfpw6[5] & Tfjiu6);
assign F23ju6 = (Cyfpw6[0] & Hs0iu6);
assign Prcpw6 = (Wrcpw6 & Obbow6);
assign Obbow6 = (~(Jcaiu6 | Mr0iu6));
assign Wrcpw6 = (Dscpw6 & Lkaiu6);
assign Lkaiu6 = (!Gwyiu6);
assign Gwyiu6 = (Cyfpw6[5] & Ii0iu6);
assign Dscpw6 = (U4kiu6 | Buaow6);
assign Buaow6 = (Tr0iu6 & Xe8iu6);
assign Brcpw6 = (Kscpw6 & Rscpw6);
assign Rscpw6 = (~(Yscpw6 & W2aow6));
assign W2aow6 = (Cyfpw6[5] & Hs0iu6);
assign Yscpw6 = (~(Mr0iu6 | Y7ghu6));
assign Kscpw6 = (~(Imaiu6 & Ftcpw6));
assign Ftcpw6 = (~(Mtcpw6 & Ttcpw6));
assign Ttcpw6 = (~(Wp0iu6 | Cyfpw6[7]));
assign Mtcpw6 = (~(Cp3ju6 | Sq3ju6));
assign Sq3ju6 = (Cyfpw6[6] & Nlaiu6);
assign Cp3ju6 = (Cyfpw6[1] & Y2oiu6);
assign Nqcpw6 = (Aucpw6 & Hucpw6);
assign Hucpw6 = (Oucpw6 & Vucpw6);
assign Vucpw6 = (~(Ae0iu6 & Cvcpw6));
assign Cvcpw6 = (~(Jvcpw6 & Qvcpw6));
assign Qvcpw6 = (~(Xvcpw6 & Pfoiu6));
assign Pfoiu6 = (Xe8iu6 & Hs0iu6);
assign Hs0iu6 = (!Cyfpw6[7]);
assign Xvcpw6 = (Frziu6 & Cyfpw6[0]);
assign Frziu6 = (~(Tfjiu6 | H4ghu6));
assign Jvcpw6 = (~(Ewcpw6 & Fd0iu6));
assign Fd0iu6 = (Cyfpw6[5] & Cyfpw6[1]);
assign Ewcpw6 = (F3aiu6 & Tfjiu6);
assign Oucpw6 = (~(V9ghu6 & Lwcpw6));
assign Lwcpw6 = (~(Erhiu6 & Swcpw6));
assign Swcpw6 = (~(Zwcpw6 & Pt2ju6));
assign Pt2ju6 = (Cyfpw6[1] & Xe8iu6);
assign Zwcpw6 = (~(Qxaiu6 | Knaiu6));
assign Qxaiu6 = (!Vo3ju6);
assign Erhiu6 = (Tq9ow6 & Gxcpw6);
assign Gxcpw6 = (~(Y8aju6 & Vj9pw6));
assign Y8aju6 = (~(Nlaiu6 | Mr0iu6));
assign Tq9ow6 = (W8oiu6 | Knaiu6);
assign W8oiu6 = (!Vj9pw6);
assign Vj9pw6 = (Sbghu6 & K9aiu6);
assign Aucpw6 = (Nxcpw6 & Uxcpw6);
assign Uxcpw6 = (~(J4aju6 & Qyniu6));
assign Qyniu6 = (~(Cyfpw6[1] | Cyfpw6[6]));
assign J4aju6 = (Bycpw6 & Omyiu6);
assign Omyiu6 = (Cyfpw6[3] & Jjhiu6);
assign Bycpw6 = (~(Cyfpw6[5] | Y7ghu6));
assign Nxcpw6 = (~(Cyfpw6[4] & Iycpw6));
assign Iycpw6 = (~(Pycpw6 & Wycpw6));
assign Wycpw6 = (Dzcpw6 & Kzcpw6);
assign Kzcpw6 = (~(Z6aiu6 | N20ju6));
assign N20ju6 = (W8aiu6 & Cyfpw6[6]);
assign Z6aiu6 = (Vo3ju6 & Pugiu6);
assign Pugiu6 = (Cyfpw6[5] & Tr0iu6);
assign Dzcpw6 = (Rzcpw6 & Yzcpw6);
assign Yzcpw6 = (~(V9ghu6 & F0dpw6));
assign F0dpw6 = (~(M0dpw6 & T0dpw6));
assign T0dpw6 = (~(A1dpw6 & Vo3ju6));
assign A1dpw6 = (~(Jcaiu6 | D7fpw6[14]));
assign Jcaiu6 = (!Llaow6);
assign M0dpw6 = (~(H1dpw6 & Mr0iu6));
assign H1dpw6 = (~(O1dpw6 & V1dpw6));
assign V1dpw6 = (~(C2dpw6 & Kxziu6));
assign Kxziu6 = (~(Ae0iu6 | D7fpw6[14]));
assign C2dpw6 = (~(Ii0iu6 | Hbbow6));
assign Hbbow6 = (Dcziu6 & J2dpw6);
assign J2dpw6 = (Dzjiu6 | A1kiu6);
assign A1kiu6 = (!D7fpw6[4]);
assign Dzjiu6 = (!D7fpw6[5]);
assign O1dpw6 = (~(Llaow6 & Q2dpw6));
assign Q2dpw6 = (~(X2dpw6 & Mpaow6));
assign Mpaow6 = (~(Y40ju6 | Vk9ow6));
assign Vk9ow6 = (X1ziu6 & Ftjiu6);
assign Y40ju6 = (D7fpw6[12] & X1ziu6);
assign X2dpw6 = (~(E3dpw6 | Jiiiu6));
assign Jiiiu6 = (Uriiu6 & Ftjiu6);
assign E3dpw6 = (Ya1ju6 & D7fpw6[14]);
assign Ya1ju6 = (~(Ftjiu6 | D7fpw6[12]));
assign Llaow6 = (~(Ae0iu6 | Y7ghu6));
assign Rzcpw6 = (~(K2aiu6 & D6kiu6));
assign D6kiu6 = (~(Tfjiu6 | K9aiu6));
assign K2aiu6 = (Ii0iu6 & Xe8iu6);
assign Pycpw6 = (~(L3dpw6 | S3dpw6));
assign S3dpw6 = (Sbghu6 ? W8aiu6 : Z3dpw6);
assign Z3dpw6 = (~(Knaiu6 | Tr0iu6));
assign L3dpw6 = (~(G4dpw6 & N4dpw6));
assign N4dpw6 = (K9bow6 | Xkaow6);
assign Xkaow6 = (!Hiaiu6);
assign Hiaiu6 = (Zraiu6 & Geaiu6);
assign K9bow6 = (!X97ow6);
assign X97ow6 = (Cyfpw6[5] & Mr0iu6);
assign G4dpw6 = (P1bow6 | Nlaiu6);
assign P1bow6 = (!Neoiu6);
assign Neoiu6 = (Cyfpw6[1] & Zraiu6);
assign Zraiu6 = (!Ae0iu6);
assign Lpcpw6 = (Sufpw6[0] | Sufpw6[1]);
assign CODEHINTDE[2] = (~(U4dpw6 & B5dpw6));
assign B5dpw6 = (I5dpw6 & P5dpw6);
assign P5dpw6 = (~(W5dpw6 | Nriiu6));
assign Nriiu6 = (D6dpw6 & Vboiu6);
assign D6dpw6 = (~(E4jiu6 | Cyfpw6[5]));
assign E4jiu6 = (!Hzziu6);
assign Hzziu6 = (Cyfpw6[4] & Jjhiu6);
assign W5dpw6 = (K6dpw6 & De6ow6);
assign De6ow6 = (~(Vwaiu6 | C0ehu6));
assign Vwaiu6 = (!Wp0iu6);
assign Wp0iu6 = (Cyfpw6[0] & Xe8iu6);
assign Xe8iu6 = (!Cyfpw6[5]);
assign K6dpw6 = (~(As0iu6 | Knaiu6));
assign As0iu6 = (!Ldoiu6);
assign Ldoiu6 = (~(Tfjiu6 | Cyfpw6[4]));
assign I5dpw6 = (R6dpw6 & Y6dpw6);
assign Y6dpw6 = (~(F7dpw6 & F3aiu6));
assign F3aiu6 = (Vo3ju6 & Mr0iu6);
assign Vo3ju6 = (~(Nlaiu6 | Ii0iu6));
assign F7dpw6 = (~(Qjaiu6 | C0ehu6));
assign Qjaiu6 = (!U4kiu6);
assign U4kiu6 = (Tr0iu6 & Y2oiu6);
assign R6dpw6 = (~(Cyfpw6[7] & M7dpw6));
assign M7dpw6 = (~(Fmjiu6 & T7dpw6));
assign T7dpw6 = (Uvziu6 | Cyfpw6[0]);
assign Uvziu6 = (!Gsbow6);
assign Gsbow6 = (Cyfpw6[3] & Y7ghu6);
assign Fmjiu6 = (~(Pthiu6 & Y7ghu6));
assign U4dpw6 = (A8dpw6 & H8dpw6);
assign H8dpw6 = (O8dpw6 & V8dpw6);
assign V8dpw6 = (~(C9dpw6 & Ii0iu6));
assign Ii0iu6 = (!Cyfpw6[3]);
assign C9dpw6 = (~(J9dpw6 & Q9dpw6));
assign Q9dpw6 = (~(W8aiu6 | Ae0iu6));
assign W8aiu6 = (Y7ghu6 & Mr0iu6);
assign J9dpw6 = (X9dpw6 & Kq0iu6);
assign Kq0iu6 = (!It2ju6);
assign It2ju6 = (Y7ghu6 & Y2oiu6);
assign Y2oiu6 = (!Cyfpw6[4]);
assign X9dpw6 = (Pd6ow6 | Sbghu6);
assign Pd6ow6 = (~(Eadpw6 & D1piu6));
assign D1piu6 = (~(Nlaiu6 | C0ehu6));
assign Eadpw6 = (~(Wfoiu6 | Knaiu6));
assign Knaiu6 = (!Oiaiu6);
assign Oiaiu6 = (Cyfpw6[7] & Mr0iu6);
assign Mr0iu6 = (!H4ghu6);
assign Wfoiu6 = (!Vboiu6);
assign Vboiu6 = (Cyfpw6[6] & Tr0iu6);
assign Tr0iu6 = (!Cyfpw6[1]);
assign O8dpw6 = (S5qow6 | Y31ju6);
assign Y31ju6 = (Q5aiu6 & Uriiu6);
assign Uriiu6 = (!S1ehu6);
assign S5qow6 = (!Imaiu6);
assign Imaiu6 = (C0ehu6 & Geaiu6);
assign A8dpw6 = (Pmbow6 & Ladpw6);
assign Ladpw6 = (~(Sadpw6 & Geaiu6));
assign Sadpw6 = (~(Zadpw6 & Gbdpw6));
assign Gbdpw6 = (Nbdpw6 & Ubdpw6);
assign Ubdpw6 = (~(Bcdpw6 & J5iow6));
assign J5iow6 = (Icdpw6 & D7fpw6[14]);
assign Icdpw6 = (~(D7fpw6[13] | D7fpw6[15]));
assign Bcdpw6 = (P0piu6 & Pcdpw6);
assign Pcdpw6 = (~(Qjiow6 & Wcdpw6));
assign Wcdpw6 = (L7aow6 | I6jiu6);
assign I6jiu6 = (!D7fpw6[10]);
assign L7aow6 = (Rg2ju6 | D7fpw6[8]);
assign Rg2ju6 = (~(Dddpw6 & Kddpw6));
assign Kddpw6 = (~(Ccaiu6 | Prjiu6));
assign Prjiu6 = (!D7fpw6[2]);
assign Dddpw6 = (~(O95iu6 | Rb8iu6));
assign Qjiow6 = (!Q6aow6);
assign Q6aow6 = (Qxoiu6 & D7fpw6[8]);
assign P0piu6 = (Mtjiu6 & Oviiu6);
assign Mtjiu6 = (C0ehu6 & Gkiiu6);
assign Gkiiu6 = (!D7fpw6[12]);
assign Nbdpw6 = (~(Rddpw6 & A95iu6));
assign A95iu6 = (~(N38ow6 | D7fpw6[10]));
assign N38ow6 = (!Xiiiu6);
assign Xiiiu6 = (D7fpw6[13] & C0ehu6);
assign Rddpw6 = (Aujiu6 & Yddpw6);
assign Yddpw6 = (~(Fedpw6 & Medpw6));
assign Medpw6 = (Kcziu6 | Oviiu6);
assign Kcziu6 = (!L01ju6);
assign L01ju6 = (D7fpw6[7] & Ad8iu6);
assign Ad8iu6 = (!D7fpw6[6]);
assign Fedpw6 = (~(Il3ju6 | D7fpw6[8]));
assign Aujiu6 = (D7fpw6[15] & D7fpw6[12]);
assign Zadpw6 = (Tedpw6 & Afdpw6);
assign Afdpw6 = (~(J9kiu6 & Hfdpw6));
assign Hfdpw6 = (~(Co6ow6 & Ofdpw6));
assign Ofdpw6 = (~(D7fpw6[12] & Vfdpw6));
assign Vfdpw6 = (~(Cgdpw6 & Jgdpw6));
assign Jgdpw6 = (~(D7fpw6[13] & Qgdpw6));
assign Qgdpw6 = (Xgdpw6 | Ehdpw6);
assign Ehdpw6 = (Lhdpw6 & Qxoiu6);
assign Lhdpw6 = (~(Cwiiu6 | D7fpw6[11]));
assign Cwiiu6 = (Dcziu6 & D7fpw6[5]);
assign Dcziu6 = (D7fpw6[6] & O95iu6);
assign Xgdpw6 = (D7fpw6[8] ? Shdpw6 : F6ziu6);
assign Shdpw6 = (~(Zhdpw6 & Gidpw6));
assign Gidpw6 = (Oviiu6 | Wh0ju6);
assign Wh0ju6 = (Nidpw6 & R9aiu6);
assign R9aiu6 = (Rb8iu6 & Ccaiu6);
assign Ccaiu6 = (!D7fpw6[1]);
assign Rb8iu6 = (!D7fpw6[0]);
assign Nidpw6 = (~(D7fpw6[2] | D7fpw6[3]));
assign Zhdpw6 = (~(Zroiu6 | Il3ju6));
assign Il3ju6 = (D7fpw6[11] & Tniiu6);
assign Tniiu6 = (!D7fpw6[9]);
assign Zroiu6 = (D7fpw6[9] & Oviiu6);
assign Cgdpw6 = (~(F6ziu6 & D7fpw6[14]));
assign F6ziu6 = (Qxoiu6 & D7fpw6[11]);
assign Co6ow6 = (!Hl8ow6);
assign Hl8ow6 = (D7fpw6[13] & D7fpw6[14]);
assign J9kiu6 = (~(Jjhiu6 | Ftjiu6));
assign Ftjiu6 = (!D7fpw6[15]);
assign Tedpw6 = (Ntgiu6 | Cyfpw6[1]);
assign Ntgiu6 = (~(Pthiu6 & Yljiu6));
assign Pthiu6 = (Nlaiu6 & Tfjiu6);
assign Tfjiu6 = (!Cyfpw6[6]);
assign Pmbow6 = (Faaiu6 & Uidpw6);
assign Uidpw6 = (~(Xmliu6 & Bjdpw6));
assign Bjdpw6 = (~(Ijdpw6 & Pjdpw6));
assign Pjdpw6 = (~(Wjdpw6 & Yljiu6));
assign Wjdpw6 = (~(Cyfpw6[1] | Cyfpw6[7]));
assign Ijdpw6 = (G7oiu6 | Iuniu6);
assign Iuniu6 = (!S6aiu6);
assign S6aiu6 = (Yljiu6 & H4ghu6);
assign Yljiu6 = (Jjhiu6 & K9aiu6);
assign G7oiu6 = (!L78ju6);
assign L78ju6 = (Cyfpw6[4] & Nlaiu6);
assign Nlaiu6 = (!Cyfpw6[0]);
assign Xmliu6 = (!Taaiu6);
assign Taaiu6 = (~(Dkdpw6 & Kkdpw6));
assign Kkdpw6 = (Rkdpw6 & vis_pc_o[27]);
assign Rkdpw6 = (~(Noliu6 | Hlliu6));
assign Hlliu6 = (Ykdpw6 & H9row6);
assign H9row6 = (~(vis_ipsr_o[4] | vis_ipsr_o[5]));
assign Ykdpw6 = (Ukbpw6 & M8row6);
assign M8row6 = (~(vis_ipsr_o[2] | vis_ipsr_o[3]));
assign Ukbpw6 = (~(vis_ipsr_o[0] | vis_ipsr_o[1]));
assign Noliu6 = (!T6ehu6);
assign Dkdpw6 = (Fldpw6 & vis_pc_o[30]);
assign Fldpw6 = (vis_pc_o[29] & vis_pc_o[28]);
assign Faaiu6 = (!O4oiu6);
assign O4oiu6 = (Ae0iu6 & K9aiu6);
assign K9aiu6 = (!Y7ghu6);
assign CODEHINTDE[1] = (~(Oi2ju6 | O95iu6));
assign O95iu6 = (!D7fpw6[7]);
assign CODEHINTDE[0] = (~(Oi2ju6 | D7fpw6[7]));
assign Oi2ju6 = (!Wf2ju6);
assign Wf2ju6 = (Mldpw6 & Tldpw6);
assign Tldpw6 = (Amdpw6 & Geaiu6);
assign Geaiu6 = (!Sbghu6);
assign Amdpw6 = (Uyiiu6 | Hmdpw6);
assign Hmdpw6 = (~(Lraiu6 | Qxoiu6));
assign Qxoiu6 = (D7fpw6[10] & D7fpw6[9]);
assign Uyiiu6 = (Q5aiu6 & Oviiu6);
assign Oviiu6 = (!D7fpw6[11]);
assign Q5aiu6 = (!Lraiu6);
assign Lraiu6 = (Pzwiu6 & Cqaiu6);
assign Cqaiu6 = (!E6phu6);
assign Pzwiu6 = (Vchhu6 & Jehhu6);
assign Mldpw6 = (R7jiu6 & Ia8iu6);
assign Ia8iu6 = (~(X1ziu6 | Ae0iu6));
assign Ae0iu6 = (~(Vncpw6 | E6phu6));
assign Vncpw6 = (!Fvdhu6);
assign X1ziu6 = (!D7fpw6[14]);
assign R7jiu6 = (Ozziu6 & D7fpw6[15]);
assign Ozziu6 = (Nbkiu6 & D7fpw6[12]);
assign Nbkiu6 = (~(Jjhiu6 | D7fpw6[13]));
assign Jjhiu6 = (!C0ehu6);

always @(posedge SWCLKTCK or negedge PORESETn)
  if(~PORESETn)
    Evhpw6 <= 1'b0;
  else
    Evhpw6 <= 1'b1;

always @(posedge SWCLKTCK or negedge PORESETn)
  if(~PORESETn)
    Hwhpw6 <= 1'b0;
  else
    Hwhpw6 <= Qmdhu6;

always @(posedge SWCLKTCK or negedge PORESETn)
  if(~PORESETn)
    Kxhpw6 <= 1'b0;
  else
    Kxhpw6 <= Pndhu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Nyhpw6 <= 1'b0;
  else
    Nyhpw6 <= CDBGPWRUPACK;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    T0ipw6 <= 1'b0;
  else
    T0ipw6 <= O5ohu6;

always @(posedge DCLK) A3ipw6 <= X3yhu6;
always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    A5ipw6 <= 1'b0;
  else
    A5ipw6 <= Nrxhu6;

always @(posedge SWCLKTCK) W6ipw6 <= Grxhu6;
always @(posedge SWCLKTCK) M8ipw6 <= Jpxhu6;
always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Qaipw6 <= 1'b0;
  else
    Qaipw6 <= Sgthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Tcipw6 <= 1'b0;
  else
    Tcipw6 <= Jyohu6;

always @(posedge HCLK) Weipw6 <= Vcvhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Wgipw6 <= 1'b0;
  else
    Wgipw6 <= Fkthu6;

always @(posedge SCLK) Xiipw6 <= U1vhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Wkipw6 <= 1'b1;
  else
    Wkipw6 <= Bithu6;

always @(posedge HCLK) Vmipw6 <= Vxohu6;
always @(posedge HCLK) Uoipw6 <= Wxshu6;
always @(posedge HCLK) Uqipw6 <= Oiphu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Usipw6 <= 1'b0;
  else
    Usipw6 <= Fxuhu6;

always @(posedge HCLK) Vuipw6 <= Kyshu6;
always @(posedge HCLK) Uwipw6 <= Igvhu6;
always @(posedge HCLK) Tyipw6 <= Diuhu6;
always @(posedge SCLK) V0jpw6 <= Rbuhu6;
always @(posedge HCLK) X2jpw6 <= P6rhu6;
always @(posedge HCLK) X4jpw6 <= T8rhu6;
always @(posedge HCLK) X6jpw6 <= Hkuhu6;
always @(posedge SCLK) Z8jpw6 <= N9uhu6;
always @(posedge HCLK) Bbjpw6 <= Z5qhu6;
always @(posedge HCLK) Bdjpw6 <= D8qhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Bfjpw6 <= 1'b1;
  else
    Bfjpw6 <= Ksrhu6;

always @(posedge HCLK) Vgjpw6 <= Oxohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Qijpw6 <= 1'b0;
  else
    Qijpw6 <= Bgvhu6;

always @(posedge HCLK) Kkjpw6 <= Ourhu6;
always @(posedge HCLK) Kmjpw6 <= Zwrhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Kojpw6 <= 1'b0;
  else
    Kojpw6 <= Mxuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Lqjpw6 <= 1'b1;
  else
    Lqjpw6 <= Hxohu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Isjpw6 <= 1'b0;
  else
    Isjpw6 <= E5xhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Aujpw6 <= 1'b0;
  else
    Aujpw6 <= Axohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Yvjpw6 <= 1'b0;
  else
    Yvjpw6 <= Twohu6;

always @(posedge HCLK) Wxjpw6 <= Mwohu6;
always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Vzjpw6 <= 1'b0;
  else
    Vzjpw6 <= Fivhu6;

always @(posedge HCLK) U1kpw6 <= Vethu6;
always @(posedge HCLK) T3kpw6 <= Amshu6;
always @(posedge HCLK) S5kpw6 <= Soshu6;
always @(posedge HCLK) R7kpw6 <= Kiuhu6;
always @(posedge SCLK) T9kpw6 <= Kbuhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Vbkpw6 <= 1'b0;
  else
    Vbkpw6 <= C6vhu6;

always @(posedge HCLK) Rdkpw6 <= Ebrhu6;
always @(posedge HCLK) Rfkpw6 <= Idrhu6;
always @(posedge HCLK) Rhkpw6 <= Okuhu6;
always @(posedge SCLK) Tjkpw6 <= G9uhu6;
always @(posedge HCLK) Vlkpw6 <= Oaqhu6;
always @(posedge HCLK) Vnkpw6 <= Scqhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Vpkpw6 <= 1'b0;
  else
    Vpkpw6 <= Bfphu6;

always @(posedge DCLK) Nrkpw6 <= I8phu6;
always @(posedge SWCLKTCK) Stkpw6 <= D0yhu6;
always @(posedge SWCLKTCK) Jvkpw6 <= Ejxhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Oxkpw6 <= 1'b0;
  else
    Oxkpw6 <= Dwuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Pzkpw6 <= 1'b1;
  else
    Pzkpw6 <= Nfvhu6;

always @(posedge HCLK) I1lpw6 <= Qdvhu6;
always @(posedge DCLK) H3lpw6 <= L6phu6;
always @(posedge SWCLKTCK) L5lpw6 <= Zqxhu6;
always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    B7lpw6 <= 1'b0;
  else
    B7lpw6 <= Fwohu6;

always @(posedge SWCLKTCK) Y8lpw6 <= Rfxhu6;
always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Kalpw6 <= 1'b1;
  else
    Kalpw6 <= Zehpw6[2];

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Bclpw6 <= 1'b0;
  else
    Bclpw6 <= Zehpw6[0];

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Sdlpw6 <= 1'b1;
  else
    Sdlpw6 <= Zehpw6[1];

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Jflpw6 <= 1'b0;
  else
    Jflpw6 <= Zehpw6[3];

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Ahlpw6 <= 1'b1;
  else
    Ahlpw6 <= Zehpw6[6];

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Rilpw6 <= 1'b1;
  else
    Rilpw6 <= Ovxhu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Yklpw6 <= 1'b0;
  else
    Yklpw6 <= Zehpw6[4];

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Pmlpw6 <= 1'b0;
  else
    Pmlpw6 <= Zehpw6[5];

always @(posedge SWCLKTCK) Golpw6 <= Yvohu6;
always @(posedge SWCLKTCK) Vplpw6 <= Rvohu6;
always @(posedge SWCLKTCK) Krlpw6 <= Kvohu6;
always @(posedge SWCLKTCK) Zslpw6 <= Dvohu6;
always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Oulpw6 <= 1'b0;
  else
    Oulpw6 <= Sqxhu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Kwlpw6 <= 1'b0;
  else
    Kwlpw6 <= Tgxhu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Gylpw6 <= 1'b0;
  else
    Gylpw6 <= Ktxhu6;

always @(posedge SWCLKTCK) Yzlpw6 <= C3yhu6;
always @(posedge SWCLKTCK) O1mpw6 <= Tnxhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    S3mpw6 <= 1'b0;
  else
    S3mpw6 <= Gvthu6;

always @(posedge SCLK) T5mpw6 <= Z0vhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    S7mpw6 <= 1'b1;
  else
    S7mpw6 <= Nhthu6;

always @(posedge HCLK) R9mpw6 <= L7vhu6;
always @(posedge HCLK) Qbmpw6 <= Wqshu6;
always @(posedge HCLK) Pdmpw6 <= Otshu6;
always @(posedge HCLK) Ofmpw6 <= Whuhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Qhmpw6 <= 1'b0;
  else
    Qhmpw6 <= Mrthu6;

always @(posedge HCLK) Mjmpw6 <= Wyrhu6;
always @(posedge HCLK) Mlmpw6 <= O1shu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Mnmpw6 <= 1'b0;
  else
    Mnmpw6 <= Xmthu6;

always @(posedge SCLK) Jpmpw6 <= N1vhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Irmpw6 <= 1'b1;
  else
    Irmpw6 <= Uhthu6;

always @(posedge HCLK) Htmpw6 <= Wuohu6;
always @(posedge HCLK) Gvmpw6 <= Ocvhu6;
always @(posedge HCLK) Gxmpw6 <= Gpshu6;
always @(posedge HCLK) Fzmpw6 <= Kkshu6;
always @(posedge HCLK) E1npw6 <= Gxrhu6;
always @(posedge HCLK) E3npw6 <= Ysrhu6;
always @(posedge HCLK) E5npw6 <= H9rhu6;
always @(posedge HCLK) E7npw6 <= S4rhu6;
always @(posedge HCLK) E9npw6 <= R8qhu6;
always @(posedge HCLK) Ebnpw6 <= C4qhu6;
always @(posedge HCLK) Ednpw6 <= Rgphu6;
always @(posedge HCLK) Efnpw6 <= Pxshu6;
always @(posedge HCLK) Ehnpw6 <= Cdvhu6;
always @(posedge HCLK) Ejnpw6 <= Jdvhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Elnpw6 <= 1'b0;
  else
    Elnpw6 <= Yjthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Fnnpw6 <= 1'b1;
  else
    Fnnpw6 <= Puohu6;

always @(posedge HCLK) Fpnpw6 <= Iuohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Arnpw6 <= 1'b1;
  else
    Arnpw6 <= Kgphu6;

always @(posedge HCLK) Usnpw6 <= Dgphu6;
always @(posedge DCLK) Uunpw6 <= H2yhu6;
always @(posedge SWCLKTCK) Zwnpw6 <= A2yhu6;
always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Qynpw6 <= 1'b0;
  else
    Qynpw6 <= Hvxhu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    I0opw6 <= 1'b0;
  else
    I0opw6 <= Q3yhu6;

always @(posedge SWCLKTCK) D2opw6 <= Wsxhu6;
always @(posedge SWCLKTCK) T3opw6 <= Hoxhu6;
always @(posedge HCLK) X5opw6 <= Gguhu6;
always @(posedge SCLK) Y7opw6 <= Oduhu6;
always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Z9opw6 <= 1'b0;
  else
    Z9opw6 <= J4xhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Xbopw6 <= 1'b1;
  else
    Xbopw6 <= N8vhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ydopw6 <= 1'b0;
  else
    Ydopw6 <= Buohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ufopw6 <= 1'b0;
  else
    Ufopw6 <= Utohu6;

always @(posedge HCLK) Shopw6 <= Ntohu6;
always @(posedge HCLK) Rjopw6 <= Evshu6;
always @(posedge HCLK) Qlopw6 <= Qushu6;
always @(posedge HCLK) Qnopw6 <= Jushu6;
always @(posedge HCLK) Qpopw6 <= Iqshu6;
always @(posedge HCLK) Propw6 <= Mlshu6;
always @(posedge HCLK) Otopw6 <= Iyrhu6;
always @(posedge HCLK) Ovopw6 <= Aurhu6;
always @(posedge HCLK) Oxopw6 <= Qarhu6;
always @(posedge HCLK) Ozopw6 <= B6rhu6;
always @(posedge HCLK) O1ppw6 <= Aaqhu6;
always @(posedge HCLK) O3ppw6 <= L5qhu6;
always @(posedge HCLK) O5ppw6 <= E9thu6;
always @(posedge HCLK) N7ppw6 <= Q8thu6;
always @(posedge HCLK) N9ppw6 <= J8thu6;
always @(posedge HCLK) Nbppw6 <= Krshu6;
always @(posedge HCLK) Mdppw6 <= Omshu6;
always @(posedge HCLK) Lfppw6 <= Kzrhu6;
always @(posedge HCLK) Lhppw6 <= Cvrhu6;
always @(posedge HCLK) Ljppw6 <= Sbrhu6;
always @(posedge HCLK) Llppw6 <= D7rhu6;
always @(posedge HCLK) Lnppw6 <= Cbqhu6;
always @(posedge HCLK) Lpppw6 <= N6qhu6;
always @(posedge HCLK) Lrppw6 <= Zevhu6;
always @(posedge HCLK) Ktppw6 <= Npshu6;
always @(posedge HCLK) Jvppw6 <= Rkshu6;
always @(posedge HCLK) Ixppw6 <= Nxrhu6;
always @(posedge HCLK) Izppw6 <= Ftrhu6;
always @(posedge HCLK) I1qpw6 <= O9rhu6;
always @(posedge HCLK) I3qpw6 <= Z4rhu6;
always @(posedge HCLK) I5qpw6 <= Y8qhu6;
always @(posedge HCLK) I7qpw6 <= J4qhu6;
always @(posedge HCLK) I9qpw6 <= Ygphu6;
always @(posedge HCLK) Ibqpw6 <= Zkphu6;
always @(posedge DCLK) Idqpw6 <= G7phu6;
always @(posedge SWCLKTCK) Nfqpw6 <= F1yhu6;
always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Ehqpw6 <= 1'b0;
  else
    Ehqpw6 <= Fgxhu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Cjqpw6 <= 1'b0;
  else
    Cjqpw6 <= Yfxhu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Xkqpw6 <= 1'b0;
  else
    Xkqpw6 <= Ytxhu6;

always @(posedge SWCLKTCK) Gnqpw6 <= Ahxhu6;
always @(posedge SWCLKTCK) Gpqpw6 <= Qpxhu6;
always @(posedge SWCLKTCK) Nrqpw6 <= Eqxhu6;
always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Utqpw6 <= 1'b0;
  else
    Utqpw6 <= Fuxhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Xvqpw6 <= 1'b0;
  else
    Xvqpw6 <= G2ohu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Xxqpw6 <= 1'b0;
  else
    Xxqpw6 <= Q7ohu6;

always @(posedge SWCLKTCK) Yzqpw6 <= V2yhu6;
always @(posedge SWCLKTCK) D2rpw6 <= Cixhu6;
always @(posedge SWCLKTCK) I4rpw6 <= Hhxhu6;
always @(posedge HCLK) M6rpw6 <= Jluhu6;
always @(posedge SCLK) N8rpw6 <= Xeuhu6;
always @(posedge SCLK) Oarpw6 <= Qeuhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Pcrpw6 <= 1'b1;
  else
    Pcrpw6 <= S0vhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Lerpw6 <= 1'b1;
  else
    Lerpw6 <= Gtohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Hgrpw6 <= 1'b1;
  else
    Hgrpw6 <= X4xhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Hirpw6 <= 1'b0;
  else
    Hirpw6 <= Zsohu6;

always @(posedge HCLK) Fkrpw6 <= Ssohu6;
always @(posedge HCLK) Emrpw6 <= Gbshu6;
always @(posedge HCLK) Dorpw6 <= Nbshu6;
always @(posedge HCLK) Cqrpw6 <= Icshu6;
always @(posedge HCLK) Bsrpw6 <= Wcshu6;
always @(posedge HCLK) Aurpw6 <= Kdshu6;
always @(posedge HCLK) Zvrpw6 <= Ofshu6;
always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Yxrpw6 <= 1'b0;
  else
    Yxrpw6 <= W1phu6;

always @(posedge HCLK) B0spw6 <= Vfshu6;
always @(posedge HCLK) A2spw6 <= Cgshu6;
always @(posedge HCLK) Z3spw6 <= Xgshu6;
always @(posedge HCLK) Y5spw6 <= Lhshu6;
always @(posedge HCLK) X7spw6 <= Zhshu6;
always @(posedge HCLK) W9spw6 <= Dkshu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Vbspw6 <= 1'b0;
  else
    Vbspw6 <= Zuthu6;

always @(posedge SCLK) Xdspw6 <= O5vhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Wfspw6 <= 1'b1;
  else
    Wfspw6 <= S7vhu6;

always @(posedge HCLK) Vhspw6 <= Lsohu6;
always @(posedge HCLK) Ujspw6 <= Fjuhu6;
always @(posedge SCLK) Wlspw6 <= Pauhu6;
always @(posedge HCLK) Ynspw6 <= K6shu6;
always @(posedge HCLK) Ypspw6 <= R6shu6;
always @(posedge HCLK) Yrspw6 <= M7shu6;
always @(posedge HCLK) Ytspw6 <= A8shu6;
always @(posedge HCLK) Yvspw6 <= O8shu6;
always @(posedge HCLK) Yxspw6 <= Sashu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Yzspw6 <= 1'b0;
  else
    Yzspw6 <= Tivhu6;

always @(posedge HCLK) Z1tpw6 <= Sirhu6;
always @(posedge HCLK) Z3tpw6 <= Zirhu6;
always @(posedge HCLK) Z5tpw6 <= Bkrhu6;
always @(posedge HCLK) Z7tpw6 <= Pkrhu6;
always @(posedge HCLK) Z9tpw6 <= Dlrhu6;
always @(posedge HCLK) Zbtpw6 <= Tmrhu6;
always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Zdtpw6 <= 1'b0;
  else
    Zdtpw6 <= Qmthu6;

always @(posedge HCLK) Yftpw6 <= Lvshu6;
always @(posedge HCLK) Xhtpw6 <= Ryshu6;
always @(posedge HCLK) Wjtpw6 <= L9thu6;
always @(posedge HCLK) Vltpw6 <= B9vhu6;
always @(posedge HCLK) Untpw6 <= I9vhu6;
always @(posedge HCLK) Tptpw6 <= Phuhu6;
always @(posedge SCLK) Vrtpw6 <= Fcuhu6;
always @(posedge HCLK) Xttpw6 <= V1shu6;
always @(posedge HCLK) Xvtpw6 <= C2shu6;
always @(posedge HCLK) Xxtpw6 <= X2shu6;
always @(posedge HCLK) Xztpw6 <= L3shu6;
always @(posedge HCLK) X1upw6 <= Z3shu6;
always @(posedge HCLK) X3upw6 <= D6shu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    X5upw6 <= 1'b0;
  else
    X5upw6 <= Rwuhu6;

always @(posedge HCLK) Y7upw6 <= Zqqhu6;
always @(posedge HCLK) Y9upw6 <= Grqhu6;
always @(posedge HCLK) Ybupw6 <= Isqhu6;
always @(posedge HCLK) Ydupw6 <= Wsqhu6;
always @(posedge HCLK) Yfupw6 <= Ktqhu6;
always @(posedge HCLK) Yhupw6 <= Avqhu6;
always @(posedge HCLK) Yjupw6 <= Mjuhu6;
always @(posedge SCLK) Amupw6 <= Iauhu6;
always @(posedge SCLK) Coupw6 <= S8uhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Equpw6 <= 1'b1;
  else
    Equpw6 <= Esohu6;

always @(posedge HCLK) Asupw6 <= Hfshu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ztupw6 <= 1'b0;
  else
    Ztupw6 <= Fbvhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Awupw6 <= 1'b1;
  else
    Awupw6 <= Xrohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Xxupw6 <= 1'b0;
  else
    Xxupw6 <= Qrohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Vzupw6 <= 1'b0;
  else
    Vzupw6 <= Jrohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    T1vpw6 <= 1'b0;
  else
    T1vpw6 <= Crohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    R3vpw6 <= 1'b0;
  else
    R3vpw6 <= Vqohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    P5vpw6 <= 1'b1;
  else
    P5vpw6 <= Oqohu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    K7vpw6 <= 1'b1;
  else
    K7vpw6 <= Vyuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    F9vpw6 <= 1'b0;
  else
    F9vpw6 <= Hqohu6;

always @(posedge DCLK) Gbvpw6 <= R9phu6;
always @(posedge SWCLKTCK) Ldvpw6 <= Uyxhu6;
always @(posedge SWCLKTCK) Cfvpw6 <= Nkxhu6;
always @(posedge HCLK) Hhvpw6 <= Akuhu6;
always @(posedge HCLK) Jjvpw6 <= D0rhu6;
always @(posedge HCLK) Jlvpw6 <= K0rhu6;
always @(posedge HCLK) Jnvpw6 <= M1rhu6;
always @(posedge HCLK) Jpvpw6 <= A2rhu6;
always @(posedge HCLK) Jrvpw6 <= O2rhu6;
always @(posedge HCLK) Jtvpw6 <= E4rhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Jvvpw6 <= 1'b0;
  else
    Jvvpw6 <= Dhvhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Dxvpw6 <= 1'b1;
  else
    Dxvpw6 <= Gfvhu6;

always @(posedge HCLK) Dzvpw6 <= Aqohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    C1wpw6 <= 1'b0;
  else
    C1wpw6 <= Hyuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    C3wpw6 <= 1'b0;
  else
    C3wpw6 <= Tbvhu6;

always @(posedge HCLK) C5wpw6 <= Kmqhu6;
always @(posedge HCLK) C7wpw6 <= Rmqhu6;
always @(posedge HCLK) C9wpw6 <= Tnqhu6;
always @(posedge HCLK) Cbwpw6 <= Hoqhu6;
always @(posedge HCLK) Cdwpw6 <= Voqhu6;
always @(posedge HCLK) Cfwpw6 <= Lqqhu6;
always @(posedge HCLK) Chwpw6 <= Sqqhu6;
always @(posedge DCLK) Cjwpw6 <= Maphu6;
always @(posedge SWCLKTCK) Hlwpw6 <= Zxxhu6;
always @(posedge SWCLKTCK) Ymwpw6 <= Ilxhu6;
always @(posedge DCLK) Dpwpw6 <= Zcxhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Sqwpw6 <= 1'b0;
  else
    Sqwpw6 <= O3xhu6;

always @(posedge DCLK) Kswpw6 <= Y9phu6;
always @(posedge SWCLKTCK) Puwpw6 <= Nyxhu6;
always @(posedge SWCLKTCK) Gwwpw6 <= Ukxhu6;
always @(posedge HCLK) Lywpw6 <= Tjuhu6;
always @(posedge SCLK) N0xpw6 <= Bauhu6;
always @(posedge HCLK) P2xpw6 <= Ovqhu6;
always @(posedge HCLK) P4xpw6 <= Vvqhu6;
always @(posedge HCLK) P6xpw6 <= Xwqhu6;
always @(posedge HCLK) P8xpw6 <= Lxqhu6;
always @(posedge HCLK) Paxpw6 <= Zxqhu6;
always @(posedge HCLK) Pcxpw6 <= Pzqhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Pexpw6 <= 1'b0;
  else
    Pexpw6 <= Khvhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Jgxpw6 <= 1'b1;
  else
    Jgxpw6 <= Iithu6;

always @(posedge HCLK) Iixpw6 <= Q4xhu6;
always @(posedge HCLK) Hkxpw6 <= Yuphu6;
always @(posedge HCLK) Hmxpw6 <= Fvphu6;
always @(posedge HCLK) Hoxpw6 <= Hwphu6;
always @(posedge HCLK) Hqxpw6 <= Vwphu6;
always @(posedge HCLK) Hsxpw6 <= Jxphu6;
always @(posedge HCLK) Huxpw6 <= Zyphu6;
always @(posedge HCLK) Gwxpw6 <= Gzphu6;
always @(posedge DCLK) Gyxpw6 <= Ccphu6;
always @(posedge SWCLKTCK) L0ypw6 <= Jwxhu6;
always @(posedge SWCLKTCK) C2ypw6 <= Ymxhu6;
always @(posedge DCLK) H4ypw6 <= Pexhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    W5ypw6 <= 1'b0;
  else
    W5ypw6 <= Yavhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    X7ypw6 <= 1'b0;
  else
    X7ypw6 <= L0vhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    U9ypw6 <= 1'b1;
  else
    U9ypw6 <= Rhvhu6;

always @(posedge HCLK) Ubypw6 <= Tpohu6;
always @(posedge HCLK) Tdypw6 <= Hnrhu6;
always @(posedge HCLK) Sfypw6 <= Onrhu6;
always @(posedge HCLK) Rhypw6 <= Qorhu6;
always @(posedge HCLK) Qjypw6 <= Eprhu6;
always @(posedge HCLK) Plypw6 <= Sprhu6;
always @(posedge HCLK) Onypw6 <= Uqrhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Npypw6 <= 1'b0;
  else
    Npypw6 <= Brrhu6;

always @(posedge HCLK) Jrypw6 <= P9vhu6;
always @(posedge HCLK) Ftypw6 <= P4thu6;
always @(posedge HCLK) Evypw6 <= I4thu6;
always @(posedge HCLK) Exypw6 <= B4thu6;
always @(posedge HCLK) Ezypw6 <= N3thu6;
always @(posedge HCLK) D1zpw6 <= Atshu6;
always @(posedge HCLK) C3zpw6 <= Eoshu6;
always @(posedge HCLK) B5zpw6 <= Pjshu6;
always @(posedge HCLK) A7zpw6 <= Afshu6;
always @(posedge HCLK) Z8zpw6 <= Eashu6;
always @(posedge HCLK) Zazpw6 <= P5shu6;
always @(posedge HCLK) Zczpw6 <= A1shu6;
always @(posedge HCLK) Zezpw6 <= Swrhu6;
always @(posedge HCLK) Zgzpw6 <= G3thu6;
always @(posedge HCLK) Yizpw6 <= Z2thu6;
always @(posedge HCLK) Ykzpw6 <= S2thu6;
always @(posedge HCLK) Ymzpw6 <= E2thu6;
always @(posedge HCLK) Xozpw6 <= Tsshu6;
always @(posedge HCLK) Wqzpw6 <= Xnshu6;
always @(posedge HCLK) Vszpw6 <= Ijshu6;
always @(posedge HCLK) Uuzpw6 <= Teshu6;
always @(posedge HCLK) Twzpw6 <= X9shu6;
always @(posedge HCLK) Tyzpw6 <= I5shu6;
always @(posedge HCLK) T00qw6 <= T0shu6;
always @(posedge HCLK) T20qw6 <= Lwrhu6;
always @(posedge HCLK) T40qw6 <= Mmrhu6;
always @(posedge HCLK) T60qw6 <= Bdrhu6;
always @(posedge HCLK) T80qw6 <= M8rhu6;
always @(posedge HCLK) Ta0qw6 <= X3rhu6;
always @(posedge HCLK) Tc0qw6 <= Izqhu6;
always @(posedge HCLK) Te0qw6 <= Tuqhu6;
always @(posedge HCLK) Tg0qw6 <= Eqqhu6;
always @(posedge HCLK) Ti0qw6 <= Lcqhu6;
always @(posedge HCLK) Tk0qw6 <= W7qhu6;
always @(posedge HCLK) Tm0qw6 <= Syphu6;
always @(posedge HCLK) So0qw6 <= Hpphu6;
always @(posedge HCLK) Rq0qw6 <= Bhuhu6;
always @(posedge SCLK) Ss0qw6 <= Tcuhu6;
always @(posedge HCLK) Tu0qw6 <= Nlphu6;
always @(posedge HCLK) Sw0qw6 <= Ulphu6;
always @(posedge HCLK) Ry0qw6 <= Wmphu6;
always @(posedge HCLK) Q01qw6 <= Knphu6;
always @(posedge HCLK) P21qw6 <= Ynphu6;
always @(posedge HCLK) O41qw6 <= Opphu6;
always @(posedge HCLK) N61qw6 <= Vpphu6;
always @(posedge DCLK) M81qw6 <= Qcphu6;
always @(posedge SWCLKTCK) Qa1qw6 <= Vvxhu6;
always @(posedge SWCLKTCK) Gc1qw6 <= Mnxhu6;
always @(posedge DCLK) Ke1qw6 <= U6xhu6;
always @(posedge DCLK) Yf1qw6 <= N6xhu6;
always @(posedge DCLK) Mh1qw6 <= Jcphu6;
always @(posedge SWCLKTCK) Qj1qw6 <= Cwxhu6;
always @(posedge SWCLKTCK) Gl1qw6 <= Fnxhu6;
always @(posedge HCLK) Kn1qw6 <= Kuphu6;
always @(posedge HCLK) Jp1qw6 <= Cqphu6;
always @(posedge HCLK) Ir1qw6 <= Jqphu6;
always @(posedge HCLK) Ht1qw6 <= Lrphu6;
always @(posedge HCLK) Gv1qw6 <= Zrphu6;
always @(posedge HCLK) Fx1qw6 <= Nsphu6;
always @(posedge HCLK) Ez1qw6 <= Btphu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    D12qw6 <= 1'b1;
  else
    D12qw6 <= Mpohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    A32qw6 <= 1'b1;
  else
    A32qw6 <= Fpohu6;

always @(posedge DCLK) X42qw6 <= S6phu6;
always @(posedge SWCLKTCK) C72qw6 <= T1yhu6;
always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    T82qw6 <= 1'b0;
  else
    T82qw6 <= Lqxhu6;

always @(posedge SWCLKTCK) Ra2qw6 <= Ohxhu6;
always @(posedge DCLK) Wc2qw6 <= F9xhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Le2qw6 <= 1'b0;
  else
    Le2qw6 <= F2xhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Dg2qw6 <= 1'b0;
  else
    Dg2qw6 <= G6xhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Uh2qw6 <= 1'b0;
  else
    Uh2qw6 <= Ghthu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Nj2qw6 <= 1'b1;
  else
    Nj2qw6 <= E7vhu6;

always @(posedge DCLK) Fl2qw6 <= B8phu6;
always @(posedge SWCLKTCK) Kn2qw6 <= K0yhu6;
always @(posedge SWCLKTCK) Bp2qw6 <= Xixhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Gr2qw6 <= 1'b0;
  else
    Gr2qw6 <= W0xhu6;

always @(posedge DCLK) Bt2qw6 <= I0xhu6;
always @(posedge DCLK) Xu2qw6 <= Zdphu6;
always @(posedge SWCLKTCK) Bx2qw6 <= Bsxhu6;
always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Ry2qw6 <= 1'b0;
  else
    Ry2qw6 <= J3yhu6;

always @(posedge SWCLKTCK) L03qw6 <= Voxhu6;
always @(posedge DCLK) P23qw6 <= D8xhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    D43qw6 <= 1'b0;
  else
    D43qw6 <= T2xhu6;

always @(posedge DCLK) V53qw6 <= Sdphu6;
always @(posedge SWCLKTCK) Z73qw6 <= Psxhu6;
always @(posedge SWCLKTCK) P93qw6 <= Ooxhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Tb3qw6 <= 1'b0;
  else
    Tb3qw6 <= Dfxhu6;

always @(posedge DCLK) Nd3qw6 <= B7xhu6;
always @(posedge DCLK) Bf3qw6 <= P7xhu6;
always @(posedge DCLK) Pg3qw6 <= W7xhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Di3qw6 <= 1'b0;
  else
    Di3qw6 <= A3xhu6;

always @(posedge DCLK) Vj3qw6 <= R8xhu6;
always @(posedge DCLK) Jl3qw6 <= Lcxhu6;
always @(posedge DCLK) Ym3qw6 <= Ecxhu6;
always @(posedge DCLK) No3qw6 <= Vaxhu6;
always @(posedge DCLK) Cq3qw6 <= M9xhu6;
always @(posedge DCLK) Rr3qw6 <= Z6phu6;
always @(posedge SWCLKTCK) Wt3qw6 <= M1yhu6;
always @(posedge SWCLKTCK) Nv3qw6 <= Vhxhu6;
always @(posedge HCLK) Sx3qw6 <= Ufvhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Sz3qw6 <= 1'b1;
  else
    Sz3qw6 <= Yoohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    P14qw6 <= 1'b1;
  else
    P14qw6 <= Wgvhu6;

always @(posedge HCLK) P34qw6 <= Xushu6;
always @(posedge HCLK) P54qw6 <= Dyshu6;
always @(posedge HCLK) Gp6ax6 <= L2thu6;
always @(posedge HCLK) Gr6ax6 <= U3thu6;
always @(posedge HCLK) Gt6ax6 <= X8thu6;
always @(posedge HCLK) Gv6ax6 <= W9vhu6;
always @(posedge HCLK) Gx6ax6 <= Davhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Gz6ax6 <= 1'b0;
  else
    Gz6ax6 <= Mkthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    F17ax6 <= 1'b0;
  else
    F17ax6 <= Rjthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    C37ax6 <= 1'b1;
  else
    C37ax6 <= Roohu6;

always @(posedge HCLK) Z47ax6 <= Dmqhu6;
always @(posedge DCLK) Z67ax6 <= Taphu6;
always @(posedge SWCLKTCK) E97ax6 <= Sxxhu6;
always @(posedge SWCLKTCK) Va7ax6 <= Plxhu6;
always @(posedge DCLK) Ad7ax6 <= Gdxhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Pe7ax6 <= 1'b0;
  else
    Pe7ax6 <= M2xhu6;

always @(posedge DCLK) Hg7ax6 <= Gephu6;
always @(posedge SWCLKTCK) Li7ax6 <= Urxhu6;
always @(posedge SWCLKTCK) Bk7ax6 <= Cpxhu6;
always @(posedge DCLK) Fm7ax6 <= P0xhu6;
always @(posedge DCLK) Xn7ax6 <= K8xhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Lp7ax6 <= 1'b0;
  else
    Lp7ax6 <= Xluhu6;

always @(posedge SCLK) Nr7ax6 <= U9uhu6;
always @(posedge SCLK) Pt7ax6 <= Ybuhu6;
always @(posedge SCLK) Rv7ax6 <= Hduhu6;
always @(posedge HCLK) Sx7ax6 <= Gdqhu6;
always @(posedge HCLK) Sz7ax6 <= Ndqhu6;
always @(posedge HCLK) S18ax6 <= Peqhu6;
always @(posedge HCLK) S38ax6 <= Dfqhu6;
always @(posedge HCLK) S58ax6 <= Rfqhu6;
always @(posedge HCLK) S78ax6 <= Ahqhu6;
always @(posedge HCLK) S98ax6 <= Hhqhu6;
always @(posedge HCLK) Sb8ax6 <= Ohqhu6;
always @(posedge DCLK) Sd8ax6 <= Abphu6;
always @(posedge SWCLKTCK) Xf8ax6 <= Lxxhu6;
always @(posedge SWCLKTCK) Oh8ax6 <= Exxhu6;
always @(posedge SWCLKTCK) Fj8ax6 <= Dmxhu6;
always @(posedge DCLK) Kl8ax6 <= Udxhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Zm8ax6 <= 1'b0;
  else
    Zm8ax6 <= H3xhu6;

always @(posedge DCLK) Ro8ax6 <= Obphu6;
always @(posedge SWCLKTCK) Wq8ax6 <= Xwxhu6;
always @(posedge SWCLKTCK) Ns8ax6 <= Kmxhu6;
always @(posedge DCLK) Su8ax6 <= Bexhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Hw8ax6 <= 1'b0;
  else
    Hw8ax6 <= Y1xhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Zx8ax6 <= 1'b0;
  else
    Zx8ax6 <= Z5xhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Vz8ax6 <= 1'b0;
  else
    Vz8ax6 <= S5xhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    R19ax6 <= 1'b0;
  else
    R19ax6 <= L5xhu6;

always @(posedge DCLK) N39ax6 <= Jrvhu6;
always @(posedge DCLK) J59ax6 <= Vqvhu6;
always @(posedge DCLK) G79ax6 <= Mpvhu6;
always @(posedge DCLK) D99ax6 <= Fpvhu6;
always @(posedge DCLK) Ab9ax6 <= Wnvhu6;
always @(posedge DCLK) Xc9ax6 <= Pnvhu6;
always @(posedge DCLK) Ue9ax6 <= Bnvhu6;
always @(posedge DCLK) Rg9ax6 <= Umvhu6;
always @(posedge DCLK) Oi9ax6 <= Gmvhu6;
always @(posedge DCLK) Lk9ax6 <= Zlvhu6;
always @(posedge DCLK) Im9ax6 <= Llvhu6;
always @(posedge DCLK) Fo9ax6 <= Xkvhu6;
always @(posedge DCLK) Bq9ax6 <= Qkvhu6;
always @(posedge DCLK) Xr9ax6 <= Ckvhu6;
always @(posedge DCLK) Tt9ax6 <= Vjvhu6;
always @(posedge DCLK) Pv9ax6 <= Ojvhu6;
always @(posedge DCLK) Lx9ax6 <= Hjvhu6;
always @(posedge DCLK) Hz9ax6 <= Ajvhu6;
always @(posedge DCLK) D1aax6 <= D2whu6;
always @(posedge DCLK) Z2aax6 <= P1whu6;
always @(posedge DCLK) W4aax6 <= G0whu6;
always @(posedge DCLK) T6aax6 <= Zzvhu6;
always @(posedge DCLK) Q8aax6 <= Qyvhu6;
always @(posedge DCLK) Naaax6 <= Jyvhu6;
always @(posedge DCLK) Kcaax6 <= Vxvhu6;
always @(posedge DCLK) Heaax6 <= Oxvhu6;
always @(posedge DCLK) Egaax6 <= Axvhu6;
always @(posedge DCLK) Biaax6 <= Twvhu6;
always @(posedge DCLK) Yjaax6 <= Fwvhu6;
always @(posedge DCLK) Vlaax6 <= Rvvhu6;
always @(posedge DCLK) Rnaax6 <= Kvvhu6;
always @(posedge DCLK) Npaax6 <= Wuvhu6;
always @(posedge DCLK) Jraax6 <= Puvhu6;
always @(posedge DCLK) Ftaax6 <= Iuvhu6;
always @(posedge DCLK) Bvaax6 <= Buvhu6;
always @(posedge DCLK) Xwaax6 <= Utvhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Tyaax6 <= 1'b0;
  else
    Tyaax6 <= Ntvhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    P0bax6 <= 1'b0;
  else
    P0bax6 <= Gtvhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    L2bax6 <= 1'b0;
  else
    L2bax6 <= Zsvhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    H4bax6 <= 1'b0;
  else
    H4bax6 <= T3whu6;

always @(posedge DCLK) X5bax6 <= Qrvhu6;
always @(posedge DCLK) T7bax6 <= Xrvhu6;
always @(posedge DCLK) P9bax6 <= Esvhu6;
always @(posedge DCLK) Lbbax6 <= Lsvhu6;
always @(posedge DCLK) Hdbax6 <= K2whu6;
always @(posedge DCLK) Dfbax6 <= R2whu6;
always @(posedge DCLK) Zgbax6 <= Y2whu6;
always @(posedge DCLK) Vibax6 <= F3whu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Rkbax6 <= 1'b0;
  else
    Rkbax6 <= Ifphu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Hmbax6 <= 1'b0;
  else
    Hmbax6 <= Oyuhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Xnbax6 <= 1'b0;
  else
    Xnbax6 <= X6vhu6;

always @(posedge DCLK) Opbax6 <= Vbwhu6;
always @(posedge DCLK) Krbax6 <= Hbwhu6;
always @(posedge DCLK) Htbax6 <= Fawhu6;
always @(posedge DCLK) Evbax6 <= Y9whu6;
always @(posedge DCLK) Bxbax6 <= P8whu6;
always @(posedge DCLK) Yybax6 <= I8whu6;
always @(posedge DCLK) V0cax6 <= U7whu6;
always @(posedge DCLK) S2cax6 <= N7whu6;
always @(posedge DCLK) P4cax6 <= Z6whu6;
always @(posedge DCLK) M6cax6 <= S6whu6;
always @(posedge DCLK) J8cax6 <= E6whu6;
always @(posedge DCLK) Facax6 <= Q5whu6;
always @(posedge DCLK) Bccax6 <= J5whu6;
always @(posedge DCLK) Xdcax6 <= V4whu6;
always @(posedge DCLK) Tfcax6 <= O4whu6;
always @(posedge DCLK) Phcax6 <= H4whu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Ljcax6 <= 1'b0;
  else
    Ljcax6 <= A4whu6;

always @(posedge DCLK) Hlcax6 <= B0xhu6;
always @(posedge DCLK) Dncax6 <= Nzwhu6;
always @(posedge DCLK) Apcax6 <= Lywhu6;
always @(posedge DCLK) Xqcax6 <= Eywhu6;
always @(posedge DCLK) Uscax6 <= Vwwhu6;
always @(posedge DCLK) Rucax6 <= Owwhu6;
always @(posedge DCLK) Owcax6 <= Awwhu6;
always @(posedge DCLK) Lycax6 <= Tvwhu6;
always @(posedge DCLK) I0dax6 <= Fvwhu6;
always @(posedge DCLK) F2dax6 <= Yuwhu6;
always @(posedge DCLK) C4dax6 <= Kuwhu6;
always @(posedge DCLK) Y5dax6 <= Wtwhu6;
always @(posedge DCLK) U7dax6 <= Ptwhu6;
always @(posedge DCLK) Q9dax6 <= Btwhu6;
always @(posedge DCLK) Mbdax6 <= Uswhu6;
always @(posedge DCLK) Iddax6 <= Nswhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Efdax6 <= 1'b0;
  else
    Efdax6 <= Gswhu6;

always @(posedge DCLK) Ahdax6 <= Zrwhu6;
always @(posedge DCLK) Widax6 <= Lrwhu6;
always @(posedge DCLK) Tkdax6 <= Jqwhu6;
always @(posedge DCLK) Qmdax6 <= Cqwhu6;
always @(posedge DCLK) Nodax6 <= Towhu6;
always @(posedge DCLK) Kqdax6 <= Mowhu6;
always @(posedge DCLK) Hsdax6 <= Ynwhu6;
always @(posedge DCLK) Eudax6 <= Rnwhu6;
always @(posedge DCLK) Bwdax6 <= Dnwhu6;
always @(posedge DCLK) Yxdax6 <= Wmwhu6;
always @(posedge DCLK) Vzdax6 <= Imwhu6;
always @(posedge DCLK) R1eax6 <= Ulwhu6;
always @(posedge DCLK) N3eax6 <= Nlwhu6;
always @(posedge DCLK) J5eax6 <= Zkwhu6;
always @(posedge DCLK) F7eax6 <= Skwhu6;
always @(posedge DCLK) B9eax6 <= Lkwhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Xaeax6 <= 1'b0;
  else
    Xaeax6 <= Ekwhu6;

always @(posedge DCLK) Tceax6 <= Xjwhu6;
always @(posedge DCLK) Peeax6 <= Jjwhu6;
always @(posedge DCLK) Mgeax6 <= Hiwhu6;
always @(posedge DCLK) Jieax6 <= Aiwhu6;
always @(posedge DCLK) Gkeax6 <= Rgwhu6;
always @(posedge DCLK) Dmeax6 <= Kgwhu6;
always @(posedge DCLK) Aoeax6 <= Wfwhu6;
always @(posedge DCLK) Xpeax6 <= Pfwhu6;
always @(posedge DCLK) Ureax6 <= Bfwhu6;
always @(posedge DCLK) Rteax6 <= Uewhu6;
always @(posedge DCLK) Oveax6 <= Gewhu6;
always @(posedge DCLK) Kxeax6 <= Sdwhu6;
always @(posedge DCLK) Gzeax6 <= Ldwhu6;
always @(posedge DCLK) C1fax6 <= Xcwhu6;
always @(posedge DCLK) Y2fax6 <= Qcwhu6;
always @(posedge DCLK) U4fax6 <= Jcwhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Q6fax6 <= 1'b0;
  else
    Q6fax6 <= Ccwhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    M8fax6 <= 1'b0;
  else
    M8fax6 <= Czuhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Eafax6 <= 1'b0;
  else
    Eafax6 <= K1xhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Sbfax6 <= 1'b0;
  else
    Sbfax6 <= R1xhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Hdfax6 <= 1'b0;
  else
    Hdfax6 <= D1xhu6;

always @(posedge DCLK) Vefax6 <= Edphu6;
always @(posedge SWCLKTCK) Zgfax6 <= Dtxhu6;
always @(posedge SWCLKTCK) Pifax6 <= Avxhu6;
always @(posedge SWCLKTCK) Okfax6 <= Isxhu6;
always @(posedge SWCLKTCK) Nmfax6 <= Xpxhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Uofax6 <= 1'b0;
  else
    Uofax6 <= Pkhpw6[1];

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Sqfax6 <= 1'b0;
  else
    Sqfax6 <= Pkhpw6[0];

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Qsfax6 <= 1'b0;
  else
    Qsfax6 <= Muxhu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Qufax6 <= 1'b0;
  else
    Qufax6 <= Dtnhu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Qwfax6 <= 1'b0;
  else
    Qwfax6 <= S3ohu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Ryfax6 <= 1'b0;
  else
    Ryfax6 <= Rtxhu6;

always @(posedge SWCLKTCK) J0gax6 <= Tuxhu6;
always @(posedge DCLK) Q2gax6 <= Crvhu6;
always @(posedge DCLK) N4gax6 <= W1whu6;
always @(posedge DCLK) K6gax6 <= Obwhu6;
always @(posedge DCLK) H8gax6 <= Qjwhu6;
always @(posedge DCLK) Eagax6 <= Srwhu6;
always @(posedge DCLK) Bcgax6 <= Uzwhu6;
always @(posedge DCLK) Ydgax6 <= O2yhu6;
always @(posedge DCLK) Nfgax6 <= Hqvhu6;
always @(posedge DCLK) Khgax6 <= B1whu6;
always @(posedge DCLK) Hjgax6 <= Abwhu6;
always @(posedge DCLK) Elgax6 <= Cjwhu6;
always @(posedge DCLK) Bngax6 <= Erwhu6;
always @(posedge DCLK) Yogax6 <= Gzwhu6;
always @(posedge DCLK) Vqgax6 <= T9xhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Ksgax6 <= 1'b0;
  else
    Ksgax6 <= Kfxhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Dugax6 <= 1'b0;
  else
    Dugax6 <= Wexhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Wvgax6 <= 1'b0;
  else
    Wvgax6 <= C4xhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Jxgax6 <= 1'b1;
  else
    Jxgax6 <= V3xhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Vygax6 <= 1'b0;
  else
    Vygax6 <= U8vhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    U0hax6 <= 1'b1;
  else
    U0hax6 <= Koohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    R2hax6 <= 1'b1;
  else
    R2hax6 <= Doohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    O4hax6 <= 1'b1;
  else
    O4hax6 <= Wnohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    L6hax6 <= 1'b1;
  else
    L6hax6 <= Pnohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    I8hax6 <= 1'b1;
  else
    I8hax6 <= Inohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Fahax6 <= 1'b1;
  else
    Fahax6 <= Bnohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Cchax6 <= 1'b1;
  else
    Cchax6 <= Umohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Zdhax6 <= 1'b1;
  else
    Zdhax6 <= Nmohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Wfhax6 <= 1'b1;
  else
    Wfhax6 <= Gmohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Thhax6 <= 1'b1;
  else
    Thhax6 <= Zlohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Qjhax6 <= 1'b1;
  else
    Qjhax6 <= Slohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Nlhax6 <= 1'b1;
  else
    Nlhax6 <= Llohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Knhax6 <= 1'b1;
  else
    Knhax6 <= Elohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Hphax6 <= 1'b1;
  else
    Hphax6 <= Xkohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Drhax6 <= 1'b1;
  else
    Drhax6 <= Qkohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Zshax6 <= 1'b1;
  else
    Zshax6 <= Jkohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Vuhax6 <= 1'b1;
  else
    Vuhax6 <= Ckohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Rwhax6 <= 1'b1;
  else
    Rwhax6 <= Vjohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Nyhax6 <= 1'b1;
  else
    Nyhax6 <= Ojohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    J0iax6 <= 1'b1;
  else
    J0iax6 <= Hjohu6;

always @(posedge SCLK) G2iax6 <= B2vhu6;
always @(posedge SCLK) F4iax6 <= I2vhu6;
always @(posedge SCLK) E6iax6 <= H5vhu6;
always @(posedge SCLK) E8iax6 <= D3vhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Daiax6 <= 1'b0;
  else
    Daiax6 <= Ajohu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Bciax6 <= 1'b0;
  else
    Bciax6 <= P2vhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Zdiax6 <= 1'b0;
  else
    Zdiax6 <= Tiohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Xfiax6 <= 1'b0;
  else
    Xfiax6 <= Xdvhu6;

always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Thiax6 <= 1'b0;
  else
    Thiax6 <= Frthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ijiax6 <= 1'b0;
  else
    Ijiax6 <= Ctthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Eliax6 <= 1'b1;
  else
    Eliax6 <= W2vhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Aniax6 <= 1'b0;
  else
    Aniax6 <= G1vhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Woiax6 <= 1'b0;
  else
    Woiax6 <= Bpthu6;

always @(posedge SCLK) Zqiax6 <= K3vhu6;
always @(posedge SCLK) Ysiax6 <= R3vhu6;
always @(posedge SCLK) Xuiax6 <= Y3vhu6;
always @(posedge SCLK) Wwiax6 <= F4vhu6;
always @(posedge SCLK) Wyiax6 <= M4vhu6;
always @(posedge SCLK) W0jax6 <= T4vhu6;
always @(posedge SCLK) W2jax6 <= A5vhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    W4jax6 <= 1'b1;
  else
    W4jax6 <= Withu6;

always @(posedge HCLK) V6jax6 <= Miohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    U8jax6 <= 1'b0;
  else
    U8jax6 <= Fiohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Tajax6 <= 1'b1;
  else
    Tajax6 <= Yhohu6;

always @(posedge HCLK) Tcjax6 <= Rhohu6;
always @(posedge HCLK) Sejax6 <= Khohu6;
always @(posedge HCLK) Sgjax6 <= Dhohu6;
always @(posedge HCLK) Sijax6 <= Wgohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Skjax6 <= 1'b1;
  else
    Skjax6 <= E0vhu6;

always @(posedge HCLK) Smjax6 <= Pgohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Sojax6 <= 1'b1;
  else
    Sojax6 <= Xzuhu6;

always @(posedge HCLK) Sqjax6 <= Igohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ssjax6 <= 1'b1;
  else
    Ssjax6 <= Qzuhu6;

always @(posedge HCLK) Sujax6 <= Bgohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Rwjax6 <= 1'b1;
  else
    Rwjax6 <= Jzuhu6;

always @(posedge HCLK) Qyjax6 <= Ufohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    P0kax6 <= 1'b1;
  else
    P0kax6 <= V5vhu6;

always @(posedge HCLK) O2kax6 <= Nfohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    N4kax6 <= 1'b1;
  else
    N4kax6 <= Djthu6;

always @(posedge HCLK) M6kax6 <= Gfohu6;
always @(posedge HCLK) L8kax6 <= Zeohu6;
always @(posedge HCLK) Kakax6 <= Seohu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Jckax6 <= 1'b1;
  else
    Jckax6 <= Pithu6;

always @(posedge HCLK) Iekax6 <= Xfthu6;
always @(posedge HCLK) Lgkax6 <= Qfthu6;
always @(posedge HCLK) Oikax6 <= Jfthu6;
always @(posedge HCLK) Rkkax6 <= Cfthu6;
always @(posedge HCLK) Umkax6 <= Leohu6;
always @(posedge HCLK) Tokax6 <= Eeohu6;
always @(posedge HCLK) Sqkax6 <= Pgvhu6;
always @(posedge HCLK) Rskax6 <= Oethu6;
always @(posedge HCLK) Qukax6 <= Cushu6;
always @(posedge HCLK) Pwkax6 <= Ixshu6;
always @(posedge HCLK) Oykax6 <= C8thu6;
always @(posedge HCLK) N0lax6 <= Eevhu6;
always @(posedge HCLK) M2lax6 <= Sevhu6;
always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    L4lax6 <= 1'b1;
  else
    L4lax6 <= Wfphu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    L6lax6 <= 1'b1;
  else
    L6lax6 <= Xdohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    I8lax6 <= 1'b0;
  else
    I8lax6 <= Qdohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Halax6 <= 1'b0;
  else
    Halax6 <= Z7vhu6;

always @(posedge HCLK) Eclax6 <= Bxshu6;
always @(posedge HCLK) Delax6 <= Uwshu6;
always @(posedge HCLK) Cglax6 <= Nwshu6;
always @(posedge HCLK) Cilax6 <= Gwshu6;
always @(posedge HCLK) Cklax6 <= Zvshu6;
always @(posedge HCLK) Cmlax6 <= Svshu6;
always @(posedge HCLK) Bolax6 <= Pqshu6;
always @(posedge HCLK) Aqlax6 <= Tlshu6;
always @(posedge HCLK) Zrlax6 <= Ehshu6;
always @(posedge HCLK) Ytlax6 <= Pcshu6;
always @(posedge HCLK) Xvlax6 <= T7shu6;
always @(posedge HCLK) Xxlax6 <= E3shu6;
always @(posedge HCLK) Xzlax6 <= Pyrhu6;
always @(posedge HCLK) X1max6 <= Hurhu6;
always @(posedge HCLK) X3max6 <= Xorhu6;
always @(posedge HCLK) W5max6 <= Ikrhu6;
always @(posedge HCLK) W7max6 <= Xarhu6;
always @(posedge HCLK) W9max6 <= I6rhu6;
always @(posedge HCLK) Wbmax6 <= T1rhu6;
always @(posedge HCLK) Wdmax6 <= Exqhu6;
always @(posedge HCLK) Wfmax6 <= Psqhu6;
always @(posedge HCLK) Whmax6 <= Aoqhu6;
always @(posedge HCLK) Wjmax6 <= Weqhu6;
always @(posedge HCLK) Wlmax6 <= Haqhu6;
always @(posedge HCLK) Wnmax6 <= S5qhu6;
always @(posedge HCLK) Wpmax6 <= Owphu6;
always @(posedge HCLK) Wrmax6 <= Srphu6;
always @(posedge HCLK) Vtmax6 <= Dnphu6;
always @(posedge HCLK) Uvmax6 <= X1thu6;
always @(posedge HCLK) Txmax6 <= Q1thu6;
always @(posedge HCLK) Szmax6 <= J1thu6;
always @(posedge HCLK) S1nax6 <= C1thu6;
always @(posedge HCLK) S3nax6 <= V0thu6;
always @(posedge HCLK) S5nax6 <= O0thu6;
always @(posedge HCLK) R7nax6 <= Msshu6;
always @(posedge HCLK) Q9nax6 <= Qnshu6;
always @(posedge HCLK) Pbnax6 <= Bjshu6;
always @(posedge HCLK) Odnax6 <= Meshu6;
always @(posedge HCLK) Nfnax6 <= Q9shu6;
always @(posedge HCLK) Nhnax6 <= B5shu6;
always @(posedge HCLK) Njnax6 <= M0shu6;
always @(posedge HCLK) Nlnax6 <= Ewrhu6;
always @(posedge HCLK) Nnnax6 <= Fmrhu6;
always @(posedge HCLK) Npnax6 <= Ucrhu6;
always @(posedge HCLK) Nrnax6 <= F8rhu6;
always @(posedge HCLK) Ntnax6 <= Q3rhu6;
always @(posedge HCLK) Nvnax6 <= Bzqhu6;
always @(posedge HCLK) Nxnax6 <= Muqhu6;
always @(posedge HCLK) Nznax6 <= Xpqhu6;
always @(posedge HCLK) N1oax6 <= Tgqhu6;
always @(posedge HCLK) N3oax6 <= Ecqhu6;
always @(posedge HCLK) N5oax6 <= P7qhu6;
always @(posedge HCLK) N7oax6 <= Lyphu6;
always @(posedge HCLK) N9oax6 <= Apphu6;
always @(posedge HCLK) Mboax6 <= V7thu6;
always @(posedge HCLK) Ldoax6 <= O7thu6;
always @(posedge HCLK) Kfoax6 <= H7thu6;
always @(posedge HCLK) Khoax6 <= A7thu6;
always @(posedge HCLK) Kjoax6 <= T6thu6;
always @(posedge HCLK) Kloax6 <= M6thu6;
always @(posedge HCLK) Jnoax6 <= Rrshu6;
always @(posedge HCLK) Ipoax6 <= Vmshu6;
always @(posedge HCLK) Hroax6 <= Gishu6;
always @(posedge HCLK) Gtoax6 <= Rdshu6;
always @(posedge HCLK) Fvoax6 <= V8shu6;
always @(posedge HCLK) Fxoax6 <= G4shu6;
always @(posedge HCLK) Fzoax6 <= Rzrhu6;
always @(posedge HCLK) F1pax6 <= Jvrhu6;
always @(posedge HCLK) F3pax6 <= Zprhu6;
always @(posedge HCLK) E5pax6 <= Klrhu6;
always @(posedge HCLK) E7pax6 <= Zbrhu6;
always @(posedge HCLK) E9pax6 <= K7rhu6;
always @(posedge HCLK) Ebpax6 <= V2rhu6;
always @(posedge HCLK) Edpax6 <= Gyqhu6;
always @(posedge HCLK) Efpax6 <= Rtqhu6;
always @(posedge HCLK) Ehpax6 <= Cpqhu6;
always @(posedge HCLK) Ejpax6 <= Yfqhu6;
always @(posedge HCLK) Elpax6 <= Jbqhu6;
always @(posedge HCLK) Enpax6 <= U6qhu6;
always @(posedge HCLK) Eppax6 <= Qxphu6;
always @(posedge HCLK) Erpax6 <= Usphu6;
always @(posedge HCLK) Dtpax6 <= Fophu6;
always @(posedge HCLK) Cvpax6 <= Hethu6;
always @(posedge HCLK) Bxpax6 <= Aethu6;
always @(posedge HCLK) Azpax6 <= Tdthu6;
always @(posedge HCLK) A1qax6 <= Mdthu6;
always @(posedge HCLK) A3qax6 <= Fdthu6;
always @(posedge HCLK) A5qax6 <= Ycthu6;
always @(posedge HCLK) Z6qax6 <= Upshu6;
always @(posedge HCLK) Y8qax6 <= Ykshu6;
always @(posedge HCLK) Xaqax6 <= Jgshu6;
always @(posedge HCLK) Wcqax6 <= Ubshu6;
always @(posedge HCLK) Veqax6 <= Y6shu6;
always @(posedge HCLK) Vgqax6 <= J2shu6;
always @(posedge HCLK) Viqax6 <= Uxrhu6;
always @(posedge HCLK) Vkqax6 <= Mtrhu6;
always @(posedge HCLK) Vmqax6 <= Vnrhu6;
always @(posedge HCLK) Uoqax6 <= Gjrhu6;
always @(posedge HCLK) Uqqax6 <= V9rhu6;
always @(posedge HCLK) Usqax6 <= G5rhu6;
always @(posedge HCLK) Uuqax6 <= R0rhu6;
always @(posedge HCLK) Uwqax6 <= Cwqhu6;
always @(posedge HCLK) Uyqax6 <= Nrqhu6;
always @(posedge HCLK) U0rax6 <= Ymqhu6;
always @(posedge HCLK) U2rax6 <= Udqhu6;
always @(posedge HCLK) U4rax6 <= F9qhu6;
always @(posedge HCLK) U6rax6 <= Q4qhu6;
always @(posedge HCLK) U8rax6 <= Mvphu6;
always @(posedge HCLK) Uarax6 <= Qqphu6;
always @(posedge HCLK) Tcrax6 <= Bmphu6;
always @(posedge HCLK) Serax6 <= Vtshu6;
always @(posedge HCLK) Rgrax6 <= Zoshu6;
always @(posedge HCLK) Qirax6 <= Zashu6;
always @(posedge HCLK) Qkrax6 <= Rsrhu6;
always @(posedge HCLK) Qmrax6 <= Wrrhu6;
always @(posedge HCLK) Qorax6 <= Prrhu6;
always @(posedge HCLK) Pqrax6 <= Jorhu6;
always @(posedge HCLK) Osrax6 <= Ujrhu6;
always @(posedge HCLK) Ourax6 <= Jarhu6;
always @(posedge HCLK) Owrax6 <= U5rhu6;
always @(posedge HCLK) Oyrax6 <= F1rhu6;
always @(posedge HCLK) O0sax6 <= Qwqhu6;
always @(posedge HCLK) O2sax6 <= Bsqhu6;
always @(posedge HCLK) O4sax6 <= Mnqhu6;
always @(posedge HCLK) O6sax6 <= Ieqhu6;
always @(posedge HCLK) O8sax6 <= T9qhu6;
always @(posedge HCLK) Oasax6 <= E5qhu6;
always @(posedge HCLK) Ocsax6 <= Awphu6;
always @(posedge HCLK) Oesax6 <= Erphu6;
always @(posedge HCLK) Ngsax6 <= Pmphu6;
always @(posedge HCLK) Misax6 <= H0thu6;
always @(posedge HCLK) Lksax6 <= A0thu6;
always @(posedge HCLK) Kmsax6 <= Tzshu6;
always @(posedge HCLK) Kosax6 <= Mzshu6;
always @(posedge HCLK) Kqsax6 <= Fzshu6;
always @(posedge HCLK) Kssax6 <= Yyshu6;
always @(posedge HCLK) Jusax6 <= Fsshu6;
always @(posedge HCLK) Iwsax6 <= Jnshu6;
always @(posedge HCLK) Hysax6 <= Uishu6;
always @(posedge HCLK) G0tax6 <= Feshu6;
always @(posedge HCLK) F2tax6 <= J9shu6;
always @(posedge HCLK) F4tax6 <= U4shu6;
always @(posedge HCLK) F6tax6 <= F0shu6;
always @(posedge HCLK) F8tax6 <= Xvrhu6;
always @(posedge HCLK) Fatax6 <= Nqrhu6;
always @(posedge HCLK) Ectax6 <= Ylrhu6;
always @(posedge HCLK) Eetax6 <= Ncrhu6;
always @(posedge HCLK) Egtax6 <= Y7rhu6;
always @(posedge HCLK) Eitax6 <= J3rhu6;
always @(posedge HCLK) Ektax6 <= Uyqhu6;
always @(posedge HCLK) Emtax6 <= Fuqhu6;
always @(posedge HCLK) Eotax6 <= Qpqhu6;
always @(posedge HCLK) Eqtax6 <= Mgqhu6;
always @(posedge HCLK) Estax6 <= Xbqhu6;
always @(posedge HCLK) Eutax6 <= I7qhu6;
always @(posedge HCLK) Ewtax6 <= Eyphu6;
always @(posedge HCLK) Eytax6 <= Tophu6;
always @(posedge HCLK) D0uax6 <= Bbthu6;
always @(posedge HCLK) C2uax6 <= Uathu6;
always @(posedge HCLK) B4uax6 <= Nathu6;
always @(posedge HCLK) B6uax6 <= Gathu6;
always @(posedge HCLK) B8uax6 <= Z9thu6;
always @(posedge HCLK) Bauax6 <= S9thu6;
always @(posedge HCLK) Acuax6 <= Drshu6;
always @(posedge HCLK) Zduax6 <= Hmshu6;
always @(posedge HCLK) Yfuax6 <= Shshu6;
always @(posedge HCLK) Xhuax6 <= Ddshu6;
always @(posedge HCLK) Wjuax6 <= H8shu6;
always @(posedge HCLK) Wluax6 <= S3shu6;
always @(posedge HCLK) Wnuax6 <= Dzrhu6;
always @(posedge HCLK) Wpuax6 <= Vurhu6;
always @(posedge HCLK) Wruax6 <= Lprhu6;
always @(posedge HCLK) Vtuax6 <= Wkrhu6;
always @(posedge HCLK) Vvuax6 <= Lbrhu6;
always @(posedge HCLK) Vxuax6 <= W6rhu6;
always @(posedge HCLK) Vzuax6 <= H2rhu6;
always @(posedge HCLK) V1vax6 <= Sxqhu6;
always @(posedge HCLK) V3vax6 <= Dtqhu6;
always @(posedge HCLK) V5vax6 <= Ooqhu6;
always @(posedge HCLK) V7vax6 <= Kfqhu6;
always @(posedge HCLK) V9vax6 <= Vaqhu6;
always @(posedge HCLK) Vbvax6 <= G6qhu6;
always @(posedge HCLK) Vdvax6 <= Cxphu6;
always @(posedge HCLK) Vfvax6 <= Gsphu6;
always @(posedge HCLK) Uhvax6 <= Rnphu6;
always @(posedge HCLK) Tjvax6 <= F6thu6;
always @(posedge HCLK) Slvax6 <= Y5thu6;
always @(posedge HCLK) Rnvax6 <= R5thu6;
always @(posedge HCLK) Rpvax6 <= K5thu6;
always @(posedge HCLK) Rrvax6 <= D5thu6;
always @(posedge HCLK) Rtvax6 <= W4thu6;
always @(posedge HCLK) Qvvax6 <= Yrshu6;
always @(posedge HCLK) Pxvax6 <= Cnshu6;
always @(posedge HCLK) Ozvax6 <= Nishu6;
always @(posedge HCLK) N1wax6 <= Ydshu6;
always @(posedge HCLK) M3wax6 <= C9shu6;
always @(posedge HCLK) M5wax6 <= N4shu6;
always @(posedge HCLK) M7wax6 <= Yzrhu6;
always @(posedge HCLK) M9wax6 <= Qvrhu6;
always @(posedge HCLK) Mbwax6 <= Gqrhu6;
always @(posedge HCLK) Ldwax6 <= Rlrhu6;
always @(posedge HCLK) Lfwax6 <= Gcrhu6;
always @(posedge HCLK) Lhwax6 <= R7rhu6;
always @(posedge HCLK) Ljwax6 <= C3rhu6;
always @(posedge HCLK) Llwax6 <= Nyqhu6;
always @(posedge HCLK) Lnwax6 <= Ytqhu6;
always @(posedge HCLK) Lpwax6 <= Jpqhu6;
always @(posedge HCLK) Lrwax6 <= Fgqhu6;
always @(posedge HCLK) Ltwax6 <= Qbqhu6;
always @(posedge HCLK) Lvwax6 <= B7qhu6;
always @(posedge HCLK) Lxwax6 <= Xxphu6;
always @(posedge HCLK) Lzwax6 <= Mophu6;
always @(posedge HCLK) K1xax6 <= Rcthu6;
always @(posedge HCLK) J3xax6 <= Kcthu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    I5xax6 <= 1'b0;
  else
    I5xax6 <= Hcvhu6;

always @(posedge HCLK) J7xax6 <= Cluhu6;
always @(posedge HCLK) L9xax6 <= Yiuhu6;
always @(posedge SCLK) Nbxax6 <= Wauhu6;
always @(posedge HCLK) Pdxax6 <= Riuhu6;
always @(posedge SCLK) Rfxax6 <= Dbuhu6;
always @(posedge HCLK) Thxax6 <= Uguhu6;
always @(posedge SCLK) Ujxax6 <= Aduhu6;
always @(posedge HCLK) Vlxax6 <= Lfuhu6;
always @(posedge HCLK) Wnxax6 <= Efuhu6;
always @(posedge HCLK) Xpxax6 <= Zcqhu6;
always @(posedge HCLK) Xrxax6 <= Egthu6;
always @(posedge HCLK) Wtxax6 <= Lgthu6;
always @(posedge HCLK) Vvxax6 <= Dcthu6;
always @(posedge HCLK) Vxxax6 <= Wbthu6;
always @(posedge HCLK) Vzxax6 <= Pbthu6;
always @(posedge HCLK) V1yax6 <= Ibthu6;
always @(posedge HCLK) U3yax6 <= Bqshu6;
always @(posedge HCLK) T5yax6 <= Htshu6;
always @(posedge HCLK) S7yax6 <= Flshu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    R9yax6 <= 1'b0;
  else
    R9yax6 <= Mbvhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Sbyax6 <= 1'b0;
  else
    Sbyax6 <= Yqthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Pdyax6 <= 1'b0;
  else
    Pdyax6 <= Npghu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Mfyax6 <= 1'b0;
  else
    Mfyax6 <= W3uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ohyax6 <= 1'b0;
  else
    Ohyax6 <= P3uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Qjyax6 <= 1'b0;
  else
    Qjyax6 <= I3uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Slyax6 <= 1'b0;
  else
    Slyax6 <= U2uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Unyax6 <= 1'b0;
  else
    Unyax6 <= N2uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Wpyax6 <= 1'b0;
  else
    Wpyax6 <= G2uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Yryax6 <= 1'b0;
  else
    Yryax6 <= Suthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Auyax6 <= 1'b0;
  else
    Auyax6 <= Euthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Cwyax6 <= 1'b0;
  else
    Cwyax6 <= Xtthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Eyyax6 <= 1'b0;
  else
    Eyyax6 <= Qtthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    G0zax6 <= 1'b0;
  else
    G0zax6 <= Vlthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    I2zax6 <= 1'b0;
  else
    I2zax6 <= Olthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    H4zax6 <= 1'b0;
  else
    H4zax6 <= S1uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    J6zax6 <= 1'b0;
  else
    J6zax6 <= L1uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    L8zax6 <= 1'b0;
  else
    L8zax6 <= E1uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Nazax6 <= 1'b0;
  else
    Nazax6 <= Q0uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Pczax6 <= 1'b0;
  else
    Pczax6 <= J0uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Rezax6 <= 1'b0;
  else
    Rezax6 <= C0uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Tgzax6 <= 1'b0;
  else
    Tgzax6 <= Ravhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Uizax6 <= 1'b0;
  else
    Uizax6 <= Txuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Vkzax6 <= 1'b0;
  else
    Vkzax6 <= Ivuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Wmzax6 <= 1'b0;
  else
    Wmzax6 <= Aruhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Xozax6 <= 1'b0;
  else
    Xozax6 <= Mquhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Yqzax6 <= 1'b0;
  else
    Yqzax6 <= Iouhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Zszax6 <= 1'b0;
  else
    Zszax6 <= Emuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Avzax6 <= 1'b0;
  else
    Avzax6 <= Qluhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Cxzax6 <= 1'b0;
  else
    Cxzax6 <= Lmuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Czzax6 <= 1'b0;
  else
    Czzax6 <= Nnuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    C10bx6 <= 1'b0;
  else
    C10bx6 <= Pouhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    C30bx6 <= 1'b0;
  else
    C30bx6 <= Wouhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    C50bx6 <= 1'b0;
  else
    C50bx6 <= Kpuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    D70bx6 <= 1'b0;
  else
    D70bx6 <= Rpuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    E90bx6 <= 1'b0;
  else
    E90bx6 <= Ypuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Fb0bx6 <= 1'b0;
  else
    Fb0bx6 <= Fquhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Gd0bx6 <= 1'b0;
  else
    Gd0bx6 <= Tquhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Hf0bx6 <= 1'b0;
  else
    Hf0bx6 <= Hruhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ih0bx6 <= 1'b0;
  else
    Ih0bx6 <= Oruhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Jj0bx6 <= 1'b0;
  else
    Jj0bx6 <= Csuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Kl0bx6 <= 1'b0;
  else
    Kl0bx6 <= Qsuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ln0bx6 <= 1'b0;
  else
    Ln0bx6 <= Etuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Mp0bx6 <= 1'b0;
  else
    Mp0bx6 <= Stuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Nr0bx6 <= 1'b0;
  else
    Nr0bx6 <= Guuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ot0bx6 <= 1'b0;
  else
    Ot0bx6 <= Wvuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Pv0bx6 <= 1'b0;
  else
    Pv0bx6 <= Kwuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Qx0bx6 <= 1'b0;
  else
    Qx0bx6 <= Ywuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Rz0bx6 <= 1'b0;
  else
    Rz0bx6 <= Ayuhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    S11bx6 <= 1'b0;
  else
    S11bx6 <= Mivhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    U31bx6 <= 1'b0;
  else
    U31bx6 <= J5phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    W51bx6 <= 1'b0;
  else
    W51bx6 <= Gothu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Z71bx6 <= 1'b0;
  else
    Z71bx6 <= R2phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Ca1bx6 <= 1'b0;
  else
    Ca1bx6 <= Snthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Fc1bx6 <= 1'b0;
  else
    Fc1bx6 <= F3phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Ie1bx6 <= 1'b0;
  else
    Ie1bx6 <= Znthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Lg1bx6 <= 1'b0;
  else
    Lg1bx6 <= Y2phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Oi1bx6 <= 1'b0;
  else
    Oi1bx6 <= Nothu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Rk1bx6 <= 1'b0;
  else
    Rk1bx6 <= K2phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Um1bx6 <= 1'b0;
  else
    Um1bx6 <= Uothu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Xo1bx6 <= 1'b0;
  else
    Xo1bx6 <= D2phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Ar1bx6 <= 1'b0;
  else
    Ar1bx6 <= Vruhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Dt1bx6 <= 1'b0;
  else
    Dt1bx6 <= I1phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Gv1bx6 <= 1'b0;
  else
    Gv1bx6 <= Zgthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Jx1bx6 <= 1'b0;
  else
    Jx1bx6 <= P1phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Mz1bx6 <= 1'b0;
  else
    Mz1bx6 <= Jsuhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    P12bx6 <= 1'b0;
  else
    P12bx6 <= B1phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    S32bx6 <= 1'b0;
  else
    S32bx6 <= Xsuhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    V52bx6 <= 1'b0;
  else
    V52bx6 <= U0phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Y72bx6 <= 1'b0;
  else
    Y72bx6 <= Cmthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Aa2bx6 <= 1'b0;
  else
    Aa2bx6 <= C5phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Cc2bx6 <= 1'b0;
  else
    Cc2bx6 <= Ltuhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Fe2bx6 <= 1'b0;
  else
    Fe2bx6 <= N0phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Ig2bx6 <= 1'b0;
  else
    Ig2bx6 <= Ztuhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Li2bx6 <= 1'b0;
  else
    Li2bx6 <= G0phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Ok2bx6 <= 1'b0;
  else
    Ok2bx6 <= Ppthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Rm2bx6 <= 1'b0;
  else
    Rm2bx6 <= Gwdpw6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Uo2bx6 <= 1'b0;
  else
    Uo2bx6 <= Pvuhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Xq2bx6 <= 1'b0;
  else
    Xq2bx6 <= Szohu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    At2bx6 <= 1'b0;
  else
    At2bx6 <= Ipthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Dv2bx6 <= 1'b0;
  else
    Dv2bx6 <= Nwdpw6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Gx2bx6 <= 1'b0;
  else
    Gx2bx6 <= Wpthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Jz2bx6 <= 1'b0;
  else
    Jz2bx6 <= Lzohu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    M13bx6 <= 1'b0;
  else
    M13bx6 <= Dqthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    P33bx6 <= 1'b0;
  else
    P33bx6 <= Ezohu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    S53bx6 <= 1'b0;
  else
    S53bx6 <= Kqthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    V73bx6 <= 1'b0;
  else
    V73bx6 <= Xyohu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Y93bx6 <= 1'b0;
  else
    Y93bx6 <= J6vhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Bc3bx6 <= 1'b0;
  else
    Bc3bx6 <= Qyohu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Ee3bx6 <= 1'b0;
  else
    Ee3bx6 <= Q6vhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Hg3bx6 <= 1'b0;
  else
    Hg3bx6 <= Cyohu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Ki3bx6 <= 1'b0;
  else
    Ki3bx6 <= Hsthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Mk3bx6 <= 1'b0;
  else
    Mk3bx6 <= A4phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Om3bx6 <= 1'b0;
  else
    Om3bx6 <= Vsthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Qo3bx6 <= 1'b0;
  else
    Qo3bx6 <= M3phu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Sq3bx6 <= 1'b0;
  else
    Sq3bx6 <= Enthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Us3bx6 <= 1'b0;
  else
    Us3bx6 <= Bxdpw6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Wu3bx6 <= 1'b0;
  else
    Wu3bx6 <= A6uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Yw3bx6 <= 1'b0;
  else
    Yw3bx6 <= T5uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Az3bx6 <= 1'b0;
  else
    Az3bx6 <= M5uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    C14bx6 <= 1'b0;
  else
    C14bx6 <= Y4uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    E34bx6 <= 1'b0;
  else
    E34bx6 <= R4uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    G54bx6 <= 1'b0;
  else
    G54bx6 <= K4uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    I74bx6 <= 1'b0;
  else
    I74bx6 <= Kxthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    K94bx6 <= 1'b0;
  else
    K94bx6 <= Dxthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Mb4bx6 <= 1'b0;
  else
    Mb4bx6 <= Wwthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Od4bx6 <= 1'b0;
  else
    Od4bx6 <= Iwthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Qf4bx6 <= 1'b0;
  else
    Qf4bx6 <= Bwthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Sh4bx6 <= 1'b0;
  else
    Sh4bx6 <= Uvthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Uj4bx6 <= 1'b0;
  else
    Uj4bx6 <= Althu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Tl4bx6 <= 1'b0;
  else
    Tl4bx6 <= Hlthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Sn4bx6 <= 1'b0;
  else
    Sn4bx6 <= E8uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Up4bx6 <= 1'b0;
  else
    Up4bx6 <= X7uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Wr4bx6 <= 1'b0;
  else
    Wr4bx6 <= Q7uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Yt4bx6 <= 1'b0;
  else
    Yt4bx6 <= C7uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Aw4bx6 <= 1'b0;
  else
    Aw4bx6 <= V6uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Cy4bx6 <= 1'b0;
  else
    Cy4bx6 <= O6uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    E05bx6 <= 1'b0;
  else
    E05bx6 <= Ozthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    G25bx6 <= 1'b0;
  else
    G25bx6 <= Hzthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    I45bx6 <= 1'b0;
  else
    I45bx6 <= Azthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    K65bx6 <= 1'b0;
  else
    K65bx6 <= Mythu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    M85bx6 <= 1'b0;
  else
    M85bx6 <= Fythu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Oa5bx6 <= 1'b0;
  else
    Oa5bx6 <= Yxthu6;

always @(posedge HCLK) Qc5bx6 <= Loshu6;
always @(posedge HCLK) Pe5bx6 <= Qgshu6;
always @(posedge HCLK) Og5bx6 <= Bcshu6;
always @(posedge HCLK) Ni5bx6 <= F7shu6;
always @(posedge HCLK) Nk5bx6 <= Q2shu6;
always @(posedge HCLK) Nm5bx6 <= Byrhu6;
always @(posedge HCLK) No5bx6 <= Ttrhu6;
always @(posedge HCLK) Nq5bx6 <= Corhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ms5bx6 <= 1'b0;
  else
    Ms5bx6 <= Lirhu6;

always @(posedge HCLK) Nu5bx6 <= Irrhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Mw5bx6 <= 1'b1;
  else
    Mw5bx6 <= Jdohu6;

always @(posedge HCLK) Jy5bx6 <= Njrhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    J06bx6 <= 1'b1;
  else
    J06bx6 <= Cdohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    F26bx6 <= 1'b1;
  else
    F26bx6 <= Ruphu6;

always @(posedge HCLK) D46bx6 <= Carhu6;
always @(posedge HCLK) D66bx6 <= N5rhu6;
always @(posedge HCLK) D86bx6 <= Y0rhu6;
always @(posedge HCLK) Da6bx6 <= Jwqhu6;
always @(posedge HCLK) Dc6bx6 <= Urqhu6;
always @(posedge HCLK) De6bx6 <= Fnqhu6;
always @(posedge HCLK) Dg6bx6 <= Beqhu6;
always @(posedge HCLK) Di6bx6 <= M9qhu6;
always @(posedge HCLK) Dk6bx6 <= X4qhu6;
always @(posedge HCLK) Dm6bx6 <= K8qhu6;
always @(posedge HCLK) Do6bx6 <= Tvphu6;
always @(posedge HCLK) Dq6bx6 <= Xqphu6;
always @(posedge HCLK) Cs6bx6 <= Imphu6;
always @(posedge DCLK) Bu6bx6 <= Vbphu6;
always @(posedge SWCLKTCK) Gw6bx6 <= Qwxhu6;
always @(posedge SWCLKTCK) Xx6bx6 <= Rmxhu6;
always @(posedge HCLK) C07bx6 <= V3qhu6;
always @(posedge HCLK) C27bx6 <= Nzphu6;
always @(posedge HCLK) C47bx6 <= Uzphu6;
always @(posedge HCLK) C67bx6 <= B0qhu6;
always @(posedge HCLK) C87bx6 <= I0qhu6;
always @(posedge HCLK) Ca7bx6 <= P0qhu6;
always @(posedge HCLK) Cc7bx6 <= W0qhu6;
always @(posedge HCLK) Ce7bx6 <= D1qhu6;
always @(posedge HCLK) Cg7bx6 <= K1qhu6;
always @(posedge HCLK) Ci7bx6 <= R1qhu6;
always @(posedge HCLK) Ck7bx6 <= Y1qhu6;
always @(posedge HCLK) Cm7bx6 <= F2qhu6;
always @(posedge HCLK) Co7bx6 <= M2qhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Cq7bx6 <= 1'b1;
  else
    Cq7bx6 <= Vcohu6;

always @(posedge HCLK) Zr7bx6 <= Vhqhu6;
always @(posedge HCLK) Zt7bx6 <= Ciqhu6;
always @(posedge HCLK) Zv7bx6 <= Jiqhu6;
always @(posedge HCLK) Zx7bx6 <= Qiqhu6;
always @(posedge HCLK) Zz7bx6 <= Xiqhu6;
always @(posedge HCLK) Z18bx6 <= Ejqhu6;
always @(posedge HCLK) Z38bx6 <= Ljqhu6;
always @(posedge HCLK) Z58bx6 <= Sjqhu6;
always @(posedge HCLK) Z78bx6 <= Zjqhu6;
always @(posedge HCLK) Z98bx6 <= Gkqhu6;
always @(posedge HCLK) Zb8bx6 <= Nkqhu6;
always @(posedge HCLK) Zd8bx6 <= Ukqhu6;
always @(posedge HCLK) Zf8bx6 <= Blqhu6;
always @(posedge HCLK) Zh8bx6 <= Ilqhu6;
always @(posedge HCLK) Zj8bx6 <= Plqhu6;
always @(posedge HCLK) Zl8bx6 <= Wlqhu6;
always @(posedge HCLK) Zn8bx6 <= T2qhu6;
always @(posedge HCLK) Zp8bx6 <= A3qhu6;
always @(posedge HCLK) Zr8bx6 <= H3qhu6;
always @(posedge HCLK) Yt8bx6 <= O3qhu6;
always @(posedge DCLK) Xv8bx6 <= Slvhu6;
always @(posedge DCLK) Ux8bx6 <= Mwvhu6;
always @(posedge DCLK) Rz8bx6 <= L6whu6;
always @(posedge DCLK) N19bx6 <= Newhu6;
always @(posedge DCLK) J39bx6 <= Pmwhu6;
always @(posedge DCLK) F59bx6 <= Ruwhu6;
always @(posedge DCLK) B79bx6 <= Iexhu6;
always @(posedge SWCLKTCK) Q89bx6 <= Aoxhu6;
always @(posedge HCLK) Ua9bx6 <= Wjshu6;
always @(posedge DCLK) Tc9bx6 <= Jkvhu6;
always @(posedge DCLK) Pe9bx6 <= Dvvhu6;
always @(posedge DCLK) Lg9bx6 <= C5whu6;
always @(posedge DCLK) Hi9bx6 <= Edwhu6;
always @(posedge DCLK) Dk9bx6 <= Glwhu6;
always @(posedge DCLK) Zl9bx6 <= Itwhu6;
always @(posedge DCLK) Vn9bx6 <= I7xhu6;
always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Jp9bx6 <= 1'b0;
  else
    Jp9bx6 <= Osthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Lr9bx6 <= 1'b0;
  else
    Lr9bx6 <= T3phu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Nt9bx6 <= 1'b0;
  else
    Nt9bx6 <= Bouhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Nv9bx6 <= 1'b0;
  else
    Nv9bx6 <= Unuhu6;

always @(posedge HCLK) Ox9bx6 <= Nguhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Pz9bx6 <= 1'b0;
  else
    Pz9bx6 <= L8uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    R1abx6 <= 1'b0;
  else
    R1abx6 <= H6uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    T3abx6 <= 1'b0;
  else
    T3abx6 <= D4uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    V5abx6 <= 1'b0;
  else
    V5abx6 <= Z1uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    X7abx6 <= 1'b0;
  else
    X7abx6 <= Vzthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Z9abx6 <= 1'b0;
  else
    Z9abx6 <= Rxthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Bcabx6 <= 1'b0;
  else
    Bcabx6 <= Nvthu6;

always @(posedge DCLK) Ceabx6 <= Ldphu6;
always @(posedge DCLK) Ggabx6 <= Hbphu6;
always @(posedge SWCLKTCK) Liabx6 <= Wlxhu6;
always @(posedge DCLK) Qkabx6 <= Nmvhu6;
always @(posedge DCLK) Nmabx6 <= Hxvhu6;
always @(posedge DCLK) Koabx6 <= G7whu6;
always @(posedge DCLK) Hqabx6 <= Ifwhu6;
always @(posedge DCLK) Esabx6 <= Knwhu6;
always @(posedge DCLK) Buabx6 <= Mvwhu6;
always @(posedge DCLK) Yvabx6 <= Ndxhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Nxabx6 <= 1'b1;
  else
    Nxabx6 <= Ocohu6;

always @(posedge SCLK) Kzabx6 <= Jeuhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    L1bbx6 <= 1'b0;
  else
    L1bbx6 <= Smuhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    L3bbx6 <= 1'b0;
  else
    L3bbx6 <= Jmthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    N5bbx6 <= 1'b0;
  else
    N5bbx6 <= V4phu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    P7bbx6 <= 1'b1;
  else
    P7bbx6 <= Hcohu6;

always @(posedge DCLK) L9bbx6 <= Nephu6;
always @(posedge HCLK) Pbbbx6 <= Hvqhu6;
always @(posedge DCLK) Pdbbx6 <= Faphu6;
always @(posedge SWCLKTCK) Ufbbx6 <= Gyxhu6;
always @(posedge SWCLKTCK) Lhbbx6 <= Blxhu6;
always @(posedge DCLK) Qjbbx6 <= Invhu6;
always @(posedge DCLK) Nlbbx6 <= Cyvhu6;
always @(posedge DCLK) Knbbx6 <= B8whu6;
always @(posedge DCLK) Hpbbx6 <= Dgwhu6;
always @(posedge DCLK) Erbbx6 <= Fowhu6;
always @(posedge DCLK) Btbbx6 <= Hwwhu6;
always @(posedge DCLK) Yubbx6 <= Scxhu6;
always @(posedge HCLK) Nwbbx6 <= Anrhu6;
always @(posedge HCLK) Nybbx6 <= H1shu6;
always @(posedge DCLK) N0cbx6 <= N7phu6;
always @(posedge SWCLKTCK) S2cbx6 <= Y0yhu6;
always @(posedge SWCLKTCK) J4cbx6 <= R0yhu6;
always @(posedge SWCLKTCK) A6cbx6 <= Qixhu6;
always @(posedge HCLK) F8cbx6 <= W5shu6;
always @(posedge DCLK) Facbx6 <= Tpvhu6;
always @(posedge DCLK) Cccbx6 <= N0whu6;
always @(posedge DCLK) Zdcbx6 <= Mawhu6;
always @(posedge DCLK) Wfcbx6 <= Oiwhu6;
always @(posedge DCLK) Thcbx6 <= Qqwhu6;
always @(posedge DCLK) Qjcbx6 <= Sywhu6;
always @(posedge DCLK) Nlcbx6 <= Haxhu6;
always @(posedge DCLK) Cncbx6 <= U7phu6;
always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Hpcbx6 <= 1'b0;
  else
    Hpcbx6 <= Mgxhu6;

always @(posedge SWCLKTCK) Drcbx6 <= Jixhu6;
always @(posedge DCLK) Itcbx6 <= Aqvhu6;
always @(posedge DCLK) Fvcbx6 <= U0whu6;
always @(posedge DCLK) Cxcbx6 <= Tawhu6;
always @(posedge DCLK) Zycbx6 <= Viwhu6;
always @(posedge DCLK) W0dbx6 <= Xqwhu6;
always @(posedge DCLK) T2dbx6 <= Zywhu6;
always @(posedge DCLK) Q4dbx6 <= Aaxhu6;
always @(posedge HCLK) F6dbx6 <= Dsrhu6;
always @(posedge DCLK) F8dbx6 <= P8phu6;
always @(posedge SWCLKTCK) Kadbx6 <= Wzxhu6;
always @(posedge SWCLKTCK) Bcdbx6 <= Pzxhu6;
always @(posedge SWCLKTCK) Sddbx6 <= Izxhu6;
always @(posedge SWCLKTCK) Jfdbx6 <= Bzxhu6;
always @(posedge SWCLKTCK) Ahdbx6 <= Gkxhu6;
always @(posedge HCLK) Fjdbx6 <= A9rhu6;
always @(posedge DCLK) Fldbx6 <= Dovhu6;
always @(posedge DCLK) Cndbx6 <= Xyvhu6;
always @(posedge DCLK) Zodbx6 <= W8whu6;
always @(posedge DCLK) Wqdbx6 <= Ygwhu6;
always @(posedge DCLK) Tsdbx6 <= Apwhu6;
always @(posedge DCLK) Qudbx6 <= Cxwhu6;
always @(posedge DCLK) Nwdbx6 <= Xbxhu6;
always @(posedge DCLK) Cydbx6 <= K9phu6;
always @(posedge SWCLKTCK) H0ebx6 <= Zjxhu6;
always @(posedge HCLK) M2ebx6 <= Pdrhu6;
always @(posedge DCLK) M4ebx6 <= Kovhu6;
always @(posedge DCLK) J6ebx6 <= Ezvhu6;
always @(posedge DCLK) G8ebx6 <= D9whu6;
always @(posedge DCLK) Daebx6 <= Fhwhu6;
always @(posedge DCLK) Acebx6 <= Hpwhu6;
always @(posedge DCLK) Xdebx6 <= Jxwhu6;
always @(posedge DCLK) Ufebx6 <= Qbxhu6;
always @(posedge DCLK) Jhebx6 <= D9phu6;
always @(posedge SWCLKTCK) Ojebx6 <= Sjxhu6;
always @(posedge HCLK) Tlebx6 <= Eirhu6;
always @(posedge HCLK) Tnebx6 <= Wdrhu6;
always @(posedge HCLK) Tpebx6 <= Derhu6;
always @(posedge HCLK) Trebx6 <= Kerhu6;
always @(posedge HCLK) Ttebx6 <= Rerhu6;
always @(posedge HCLK) Tvebx6 <= Yerhu6;
always @(posedge HCLK) Txebx6 <= Ffrhu6;
always @(posedge HCLK) Tzebx6 <= Mfrhu6;
always @(posedge HCLK) T1fbx6 <= Tfrhu6;
always @(posedge HCLK) T3fbx6 <= Agrhu6;
always @(posedge HCLK) T5fbx6 <= Hgrhu6;
always @(posedge HCLK) T7fbx6 <= Ogrhu6;
always @(posedge HCLK) T9fbx6 <= Vgrhu6;
always @(posedge HCLK) Tbfbx6 <= Chrhu6;
always @(posedge HCLK) Tdfbx6 <= Jhrhu6;
always @(posedge HCLK) Tffbx6 <= Qhrhu6;
always @(posedge HCLK) Thfbx6 <= Xhrhu6;
always @(posedge DCLK) Tjfbx6 <= Rovhu6;
always @(posedge DCLK) Qlfbx6 <= Lzvhu6;
always @(posedge DCLK) Nnfbx6 <= K9whu6;
always @(posedge DCLK) Kpfbx6 <= Mhwhu6;
always @(posedge DCLK) Hrfbx6 <= Opwhu6;
always @(posedge DCLK) Etfbx6 <= Qxwhu6;
always @(posedge DCLK) Bvfbx6 <= Jbxhu6;
always @(posedge DCLK) Qwfbx6 <= W8phu6;
always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Vyfbx6 <= 1'b0;
  else
    Vyfbx6 <= Uuuhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Y0gbx6 <= 1'b0;
  else
    Y0gbx6 <= Zzohu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    B3gbx6 <= 1'b0;
  else
    B3gbx6 <= Bvuhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    C5gbx6 <= 1'b0;
  else
    C5gbx6 <= Nuuhu6;

always @(posedge HCLK) D7gbx6 <= Vkuhu6;
always @(posedge SCLK) F9gbx6 <= Z8uhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Hbgbx6 <= 1'b0;
  else
    Hbgbx6 <= J7uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Jdgbx6 <= 1'b0;
  else
    Jdgbx6 <= F5uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Lfgbx6 <= 1'b0;
  else
    Lfgbx6 <= B3uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Nhgbx6 <= 1'b0;
  else
    Nhgbx6 <= X0uhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Pjgbx6 <= 1'b0;
  else
    Pjgbx6 <= Tythu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Rlgbx6 <= 1'b0;
  else
    Rlgbx6 <= Pwthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Tngbx6 <= 1'b0;
  else
    Tngbx6 <= Luthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Vpgbx6 <= 1'b0;
  else
    Vpgbx6 <= Tkthu6;

always @(posedge SWCLKTCK) Urgbx6 <= Ljxhu6;
always @(posedge HCLK) Ztgbx6 <= Kavhu6;
always @(posedge DCLK) Zvgbx6 <= Yovhu6;
always @(posedge DCLK) Wxgbx6 <= Szvhu6;
always @(posedge DCLK) Tzgbx6 <= R9whu6;
always @(posedge DCLK) Q1hbx6 <= Thwhu6;
always @(posedge DCLK) N3hbx6 <= Vpwhu6;
always @(posedge DCLK) K5hbx6 <= Xxwhu6;
always @(posedge DCLK) H7hbx6 <= Cbxhu6;
always @(posedge SCLK) W8hbx6 <= Yhvhu6;
always @(posedge DCLK) Wahbx6 <= Oqvhu6;
always @(posedge DCLK) Tchbx6 <= I1whu6;
always @(posedge DCLK) Qehbx6 <= Y8xhu6;
always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Eghbx6 <= 1'b0;
  else
    Eghbx6 <= Asthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Gihbx6 <= 1'b0;
  else
    Gihbx6 <= H4phu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Ikhbx6 <= 1'b0;
  else
    Ikhbx6 <= Gnuhu6;

always @(posedge HCLK) Imhbx6 <= Zfuhu6;
always @(posedge SCLK) Johbx6 <= Vduhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Kqhbx6 <= 1'b0;
  else
    Kqhbx6 <= Jtthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Kshbx6 <= 1'b0;
  else
    Kshbx6 <= Trthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Muhbx6 <= 1'b0;
  else
    Muhbx6 <= O4phu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Owhbx6 <= 1'b0;
  else
    Owhbx6 <= Zmuhu6;

always @(posedge HCLK) Oyhbx6 <= Sfuhu6;
always @(posedge SCLK) P0ibx6 <= Ceuhu6;
always @(posedge DCLK) Q2ibx6 <= Oaxhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    F4ibx6 <= 1'b0;
  else
    F4ibx6 <= Uephu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    X5ibx6 <= 1'b0;
  else
    X5ibx6 <= Glphu6;

always @(posedge HCLK) R7ibx6 <= Fhphu6;
always @(posedge HCLK) R9ibx6 <= Mhphu6;
always @(posedge HCLK) Rbibx6 <= Thphu6;
always @(posedge HCLK) Rdibx6 <= Aiphu6;
always @(posedge HCLK) Rfibx6 <= Hiphu6;
always @(posedge HCLK) Rhibx6 <= Viphu6;
always @(posedge HCLK) Rjibx6 <= Cjphu6;
always @(posedge HCLK) Rlibx6 <= Jjphu6;
always @(posedge HCLK) Rnibx6 <= Qjphu6;
always @(posedge HCLK) Rpibx6 <= Xjphu6;
always @(posedge HCLK) Rribx6 <= Ekphu6;
always @(posedge HCLK) Rtibx6 <= Skphu6;
always @(posedge HCLK) Rvibx6 <= Itphu6;
always @(posedge HCLK) Qxibx6 <= Ptphu6;
always @(posedge HCLK) Pzibx6 <= Wtphu6;
always @(posedge HCLK) O1jbx6 <= Duphu6;
always @(posedge DCLK) N3jbx6 <= Elvhu6;
always @(posedge DCLK) J5jbx6 <= Yvvhu6;
always @(posedge DCLK) F7jbx6 <= X5whu6;
always @(posedge DCLK) B9jbx6 <= Zdwhu6;
always @(posedge DCLK) Xajbx6 <= Bmwhu6;
always @(posedge DCLK) Tcjbx6 <= Duwhu6;
always @(posedge HCLK) Pejbx6 <= Lkphu6;
always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Pgjbx6 <= 1'b0;
  else
    Pgjbx6 <= Lnthu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Rijbx6 <= 1'b0;
  else
    Rijbx6 <= Uwdpw6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Tkjbx6 <= 1'b0;
  else
    Tkjbx6 <= Dpuhu6;

always @(posedge HCLK) Tmjbx6 <= Ihuhu6;
always @(posedge SCLK) Uojbx6 <= Mcuhu6;
always @(posedge HCLK) Vqjbx6 <= Acohu6;
always @(posedge HCLK) Usjbx6 <= Tbohu6;
always @(posedge HCLK) Tujbx6 <= Mbohu6;
always @(posedge HCLK) Swjbx6 <= Fbohu6;
always @(posedge HCLK) Syjbx6 <= Wzqhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    S0kbx6 <= 1'b0;
  else
    S0kbx6 <= Acvhu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    T2kbx6 <= 1'b0;
  else
    T2kbx6 <= Kjthu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    S4kbx6 <= 1'b0;
  else
    S4kbx6 <= Levhu6;

always @(posedge HCLK) T6kbx6 <= L4rhu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    T8kbx6 <= 1'b0;
  else
    T8kbx6 <= G8vhu6;

always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Qakbx6 <= 1'b0;
  else
    Qakbx6 <= Rqthu6;

always @(posedge DCLK) Nckbx6 <= Xcphu6;
always @(posedge HCLK or negedge HRESETn)
  if(~HRESETn)
    Rekbx6 <= 1'b0;
  else
    Rekbx6 <= Yaohu6;

always @(posedge HCLK) Tgkbx6 <= Lashu6;
always @(posedge DCLK) Tikbx6 <= M3whu6;
always @(posedge DCLK) Pkkbx6 <= Ssvhu6;
always @(posedge DCLK or negedge DBGRESETn)
  if(~DBGRESETn)
    Lmkbx6 <= 1'b0;
  else
    Lmkbx6 <= Pfphu6;

always @(posedge SCLK or negedge HRESETn)
  if(~HRESETn)
    Cokbx6 <= 1'b0;
  else
    Cokbx6 <= Raohu6;

always @(posedge SWCLKTCK or negedge Fmdhu6)
  if(~Fmdhu6)
    Dqkbx6 <= 1'b0;
  else
    Dqkbx6 <= I5nhu6;

endmodule

//------------------------------------------------------------------------------
// EOF
//------------------------------------------------------------------------------

