module hello(
    input clk, reset,
    output value
);

endmodule